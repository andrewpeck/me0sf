----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- ME0 Segment Finder Firmware
-- A. Peck, A. Datta, C. Grubb, J. Chismar
----------------------------------------------------------------------------------
-- Description:
----------------------------------------------------------------------------------
library ieee;
use ieee.fixed_pkg.all;

package reciprocal_pkg is
  function reciprocal (x : integer; nbits : integer) return sfixed;
  function reciprocal6 (x : integer; nbits : integer) return sfixed;
end package reciprocal_pkg;

package body reciprocal_pkg is
  --------------------------------------------------------------------------------
  -- functions
  --------------------------------------------------------------------------------

  function reciprocal (x : integer; nbits : integer) return sfixed is
  begin
    if (x<1 or x> 2047) then
      assert false report "invalid reciprocal lookup x=" & integer'image(x) severity error;
      return to_sfixed(0, 1, -nbits);
    elsif (x=1) then return to_sfixed(1.00000000000000000000, 1, -nbits);
    elsif (x=2) then return to_sfixed(0.50000000000000000000, 1, -nbits);
    elsif (x=3) then return to_sfixed(0.33333333333333331483, 1, -nbits);
    elsif (x=4) then return to_sfixed(0.25000000000000000000, 1, -nbits);
    elsif (x=5) then return to_sfixed(0.20000000000000001110, 1, -nbits);
    elsif (x=6) then return to_sfixed(0.16666666666666665741, 1, -nbits);
    elsif (x=7) then return to_sfixed(0.14285714285714284921, 1, -nbits);
    elsif (x=8) then return to_sfixed(0.12500000000000000000, 1, -nbits);
    elsif (x=9) then return to_sfixed(0.11111111111111110494, 1, -nbits);
    elsif (x=10) then return to_sfixed(0.10000000000000000555, 1, -nbits);
    elsif (x=11) then return to_sfixed(0.09090909090909091161, 1, -nbits);
    elsif (x=12) then return to_sfixed(0.08333333333333332871, 1, -nbits);
    elsif (x=13) then return to_sfixed(0.07692307692307692735, 1, -nbits);
    elsif (x=14) then return to_sfixed(0.07142857142857142461, 1, -nbits);
    elsif (x=15) then return to_sfixed(0.06666666666666666574, 1, -nbits);
    elsif (x=16) then return to_sfixed(0.06250000000000000000, 1, -nbits);
    elsif (x=17) then return to_sfixed(0.05882352941176470507, 1, -nbits);
    elsif (x=18) then return to_sfixed(0.05555555555555555247, 1, -nbits);
    elsif (x=19) then return to_sfixed(0.05263157894736841813, 1, -nbits);
    elsif (x=20) then return to_sfixed(0.05000000000000000278, 1, -nbits);
    elsif (x=21) then return to_sfixed(0.04761904761904761640, 1, -nbits);
    elsif (x=22) then return to_sfixed(0.04545454545454545581, 1, -nbits);
    elsif (x=23) then return to_sfixed(0.04347826086956521618, 1, -nbits);
    elsif (x=24) then return to_sfixed(0.04166666666666666435, 1, -nbits);
    elsif (x=25) then return to_sfixed(0.04000000000000000083, 1, -nbits);
    elsif (x=26) then return to_sfixed(0.03846153846153846367, 1, -nbits);
    elsif (x=27) then return to_sfixed(0.03703703703703703498, 1, -nbits);
    elsif (x=28) then return to_sfixed(0.03571428571428571230, 1, -nbits);
    elsif (x=29) then return to_sfixed(0.03448275862068965469, 1, -nbits);
    elsif (x=30) then return to_sfixed(0.03333333333333333287, 1, -nbits);
    elsif (x=31) then return to_sfixed(0.03225806451612903136, 1, -nbits);
    elsif (x=32) then return to_sfixed(0.03125000000000000000, 1, -nbits);
    elsif (x=33) then return to_sfixed(0.03030303030303030387, 1, -nbits);
    elsif (x=34) then return to_sfixed(0.02941176470588235253, 1, -nbits);
    elsif (x=35) then return to_sfixed(0.02857142857142857054, 1, -nbits);
    elsif (x=36) then return to_sfixed(0.02777777777777777624, 1, -nbits);
    elsif (x=37) then return to_sfixed(0.02702702702702702853, 1, -nbits);
    elsif (x=38) then return to_sfixed(0.02631578947368420907, 1, -nbits);
    elsif (x=39) then return to_sfixed(0.02564102564102564014, 1, -nbits);
    elsif (x=40) then return to_sfixed(0.02500000000000000139, 1, -nbits);
    elsif (x=41) then return to_sfixed(0.02439024390243902524, 1, -nbits);
    elsif (x=42) then return to_sfixed(0.02380952380952380820, 1, -nbits);
    elsif (x=43) then return to_sfixed(0.02325581395348837177, 1, -nbits);
    elsif (x=44) then return to_sfixed(0.02272727272727272790, 1, -nbits);
    elsif (x=45) then return to_sfixed(0.02222222222222222307, 1, -nbits);
    elsif (x=46) then return to_sfixed(0.02173913043478260809, 1, -nbits);
    elsif (x=47) then return to_sfixed(0.02127659574468085055, 1, -nbits);
    elsif (x=48) then return to_sfixed(0.02083333333333333218, 1, -nbits);
    elsif (x=49) then return to_sfixed(0.02040816326530612082, 1, -nbits);
    elsif (x=50) then return to_sfixed(0.02000000000000000042, 1, -nbits);
    elsif (x=51) then return to_sfixed(0.01960784313725490169, 1, -nbits);
    elsif (x=52) then return to_sfixed(0.01923076923076923184, 1, -nbits);
    elsif (x=53) then return to_sfixed(0.01886792452830188607, 1, -nbits);
    elsif (x=54) then return to_sfixed(0.01851851851851851749, 1, -nbits);
    elsif (x=55) then return to_sfixed(0.01818181818181818094, 1, -nbits);
    elsif (x=56) then return to_sfixed(0.01785714285714285615, 1, -nbits);
    elsif (x=57) then return to_sfixed(0.01754385964912280604, 1, -nbits);
    elsif (x=58) then return to_sfixed(0.01724137931034482735, 1, -nbits);
    elsif (x=59) then return to_sfixed(0.01694915254237288130, 1, -nbits);
    elsif (x=60) then return to_sfixed(0.01666666666666666644, 1, -nbits);
    elsif (x=61) then return to_sfixed(0.01639344262295082053, 1, -nbits);
    elsif (x=62) then return to_sfixed(0.01612903225806451568, 1, -nbits);
    elsif (x=63) then return to_sfixed(0.01587301587301587213, 1, -nbits);
    elsif (x=64) then return to_sfixed(0.01562500000000000000, 1, -nbits);
    elsif (x=65) then return to_sfixed(0.01538461538461538547, 1, -nbits);
    elsif (x=66) then return to_sfixed(0.01515151515151515194, 1, -nbits);
    elsif (x=67) then return to_sfixed(0.01492537313432835792, 1, -nbits);
    elsif (x=68) then return to_sfixed(0.01470588235294117627, 1, -nbits);
    elsif (x=69) then return to_sfixed(0.01449275362318840597, 1, -nbits);
    elsif (x=70) then return to_sfixed(0.01428571428571428527, 1, -nbits);
    elsif (x=71) then return to_sfixed(0.01408450704225352144, 1, -nbits);
    elsif (x=72) then return to_sfixed(0.01388888888888888812, 1, -nbits);
    elsif (x=73) then return to_sfixed(0.01369863013698630061, 1, -nbits);
    elsif (x=74) then return to_sfixed(0.01351351351351351426, 1, -nbits);
    elsif (x=75) then return to_sfixed(0.01333333333333333419, 1, -nbits);
    elsif (x=76) then return to_sfixed(0.01315789473684210453, 1, -nbits);
    elsif (x=77) then return to_sfixed(0.01298701298701298787, 1, -nbits);
    elsif (x=78) then return to_sfixed(0.01282051282051282007, 1, -nbits);
    elsif (x=79) then return to_sfixed(0.01265822784810126563, 1, -nbits);
    elsif (x=80) then return to_sfixed(0.01250000000000000069, 1, -nbits);
    elsif (x=81) then return to_sfixed(0.01234567901234567833, 1, -nbits);
    elsif (x=82) then return to_sfixed(0.01219512195121951262, 1, -nbits);
    elsif (x=83) then return to_sfixed(0.01204819277108433798, 1, -nbits);
    elsif (x=84) then return to_sfixed(0.01190476190476190410, 1, -nbits);
    elsif (x=85) then return to_sfixed(0.01176470588235294101, 1, -nbits);
    elsif (x=86) then return to_sfixed(0.01162790697674418589, 1, -nbits);
    elsif (x=87) then return to_sfixed(0.01149425287356321823, 1, -nbits);
    elsif (x=88) then return to_sfixed(0.01136363636363636395, 1, -nbits);
    elsif (x=89) then return to_sfixed(0.01123595505617977497, 1, -nbits);
    elsif (x=90) then return to_sfixed(0.01111111111111111154, 1, -nbits);
    elsif (x=91) then return to_sfixed(0.01098901098901098987, 1, -nbits);
    elsif (x=92) then return to_sfixed(0.01086956521739130405, 1, -nbits);
    elsif (x=93) then return to_sfixed(0.01075268817204301161, 1, -nbits);
    elsif (x=94) then return to_sfixed(0.01063829787234042527, 1, -nbits);
    elsif (x=95) then return to_sfixed(0.01052631578947368397, 1, -nbits);
    elsif (x=96) then return to_sfixed(0.01041666666666666609, 1, -nbits);
    elsif (x=97) then return to_sfixed(0.01030927835051546372, 1, -nbits);
    elsif (x=98) then return to_sfixed(0.01020408163265306041, 1, -nbits);
    elsif (x=99) then return to_sfixed(0.01010101010101010187, 1, -nbits);
    elsif (x=100) then return to_sfixed(0.01000000000000000021, 1, -nbits);
    elsif (x=101) then return to_sfixed(0.00990099009900990111, 1, -nbits);
    elsif (x=102) then return to_sfixed(0.00980392156862745084, 1, -nbits);
    elsif (x=103) then return to_sfixed(0.00970873786407766906, 1, -nbits);
    elsif (x=104) then return to_sfixed(0.00961538461538461592, 1, -nbits);
    elsif (x=105) then return to_sfixed(0.00952380952380952467, 1, -nbits);
    elsif (x=106) then return to_sfixed(0.00943396226415094304, 1, -nbits);
    elsif (x=107) then return to_sfixed(0.00934579439252336379, 1, -nbits);
    elsif (x=108) then return to_sfixed(0.00925925925925925875, 1, -nbits);
    elsif (x=109) then return to_sfixed(0.00917431192660550510, 1, -nbits);
    elsif (x=110) then return to_sfixed(0.00909090909090909047, 1, -nbits);
    elsif (x=111) then return to_sfixed(0.00900900900900900893, 1, -nbits);
    elsif (x=112) then return to_sfixed(0.00892857142857142808, 1, -nbits);
    elsif (x=113) then return to_sfixed(0.00884955752212389368, 1, -nbits);
    elsif (x=114) then return to_sfixed(0.00877192982456140302, 1, -nbits);
    elsif (x=115) then return to_sfixed(0.00869565217391304358, 1, -nbits);
    elsif (x=116) then return to_sfixed(0.00862068965517241367, 1, -nbits);
    elsif (x=117) then return to_sfixed(0.00854700854700854787, 1, -nbits);
    elsif (x=118) then return to_sfixed(0.00847457627118644065, 1, -nbits);
    elsif (x=119) then return to_sfixed(0.00840336134453781476, 1, -nbits);
    elsif (x=120) then return to_sfixed(0.00833333333333333322, 1, -nbits);
    elsif (x=121) then return to_sfixed(0.00826446280991735560, 1, -nbits);
    elsif (x=122) then return to_sfixed(0.00819672131147541026, 1, -nbits);
    elsif (x=123) then return to_sfixed(0.00813008130081300899, 1, -nbits);
    elsif (x=124) then return to_sfixed(0.00806451612903225784, 1, -nbits);
    elsif (x=125) then return to_sfixed(0.00800000000000000017, 1, -nbits);
    elsif (x=126) then return to_sfixed(0.00793650793650793607, 1, -nbits);
    elsif (x=127) then return to_sfixed(0.00787401574803149595, 1, -nbits);
    elsif (x=128) then return to_sfixed(0.00781250000000000000, 1, -nbits);
    elsif (x=129) then return to_sfixed(0.00775193798449612392, 1, -nbits);
    elsif (x=130) then return to_sfixed(0.00769230769230769273, 1, -nbits);
    elsif (x=131) then return to_sfixed(0.00763358778625954169, 1, -nbits);
    elsif (x=132) then return to_sfixed(0.00757575757575757597, 1, -nbits);
    elsif (x=133) then return to_sfixed(0.00751879699248120259, 1, -nbits);
    elsif (x=134) then return to_sfixed(0.00746268656716417896, 1, -nbits);
    elsif (x=135) then return to_sfixed(0.00740740740740740769, 1, -nbits);
    elsif (x=136) then return to_sfixed(0.00735294117647058813, 1, -nbits);
    elsif (x=137) then return to_sfixed(0.00729927007299270049, 1, -nbits);
    elsif (x=138) then return to_sfixed(0.00724637681159420299, 1, -nbits);
    elsif (x=139) then return to_sfixed(0.00719424460431654714, 1, -nbits);
    elsif (x=140) then return to_sfixed(0.00714285714285714263, 1, -nbits);
    elsif (x=141) then return to_sfixed(0.00709219858156028352, 1, -nbits);
    elsif (x=142) then return to_sfixed(0.00704225352112676072, 1, -nbits);
    elsif (x=143) then return to_sfixed(0.00699300699300699300, 1, -nbits);
    elsif (x=144) then return to_sfixed(0.00694444444444444406, 1, -nbits);
    elsif (x=145) then return to_sfixed(0.00689655172413793094, 1, -nbits);
    elsif (x=146) then return to_sfixed(0.00684931506849315030, 1, -nbits);
    elsif (x=147) then return to_sfixed(0.00680272108843537390, 1, -nbits);
    elsif (x=148) then return to_sfixed(0.00675675675675675713, 1, -nbits);
    elsif (x=149) then return to_sfixed(0.00671140939597315422, 1, -nbits);
    elsif (x=150) then return to_sfixed(0.00666666666666666709, 1, -nbits);
    elsif (x=151) then return to_sfixed(0.00662251655629139072, 1, -nbits);
    elsif (x=152) then return to_sfixed(0.00657894736842105227, 1, -nbits);
    elsif (x=153) then return to_sfixed(0.00653594771241830085, 1, -nbits);
    elsif (x=154) then return to_sfixed(0.00649350649350649393, 1, -nbits);
    elsif (x=155) then return to_sfixed(0.00645161290322580645, 1, -nbits);
    elsif (x=156) then return to_sfixed(0.00641025641025641003, 1, -nbits);
    elsif (x=157) then return to_sfixed(0.00636942675159235701, 1, -nbits);
    elsif (x=158) then return to_sfixed(0.00632911392405063281, 1, -nbits);
    elsif (x=159) then return to_sfixed(0.00628930817610062927, 1, -nbits);
    elsif (x=160) then return to_sfixed(0.00625000000000000035, 1, -nbits);
    elsif (x=161) then return to_sfixed(0.00621118012422360206, 1, -nbits);
    elsif (x=162) then return to_sfixed(0.00617283950617283916, 1, -nbits);
    elsif (x=163) then return to_sfixed(0.00613496932515337438, 1, -nbits);
    elsif (x=164) then return to_sfixed(0.00609756097560975631, 1, -nbits);
    elsif (x=165) then return to_sfixed(0.00606060606060606060, 1, -nbits);
    elsif (x=166) then return to_sfixed(0.00602409638554216899, 1, -nbits);
    elsif (x=167) then return to_sfixed(0.00598802395209580875, 1, -nbits);
    elsif (x=168) then return to_sfixed(0.00595238095238095205, 1, -nbits);
    elsif (x=169) then return to_sfixed(0.00591715976331360933, 1, -nbits);
    elsif (x=170) then return to_sfixed(0.00588235294117647051, 1, -nbits);
    elsif (x=171) then return to_sfixed(0.00584795321637426868, 1, -nbits);
    elsif (x=172) then return to_sfixed(0.00581395348837209294, 1, -nbits);
    elsif (x=173) then return to_sfixed(0.00578034682080924827, 1, -nbits);
    elsif (x=174) then return to_sfixed(0.00574712643678160912, 1, -nbits);
    elsif (x=175) then return to_sfixed(0.00571428571428571428, 1, -nbits);
    elsif (x=176) then return to_sfixed(0.00568181818181818198, 1, -nbits);
    elsif (x=177) then return to_sfixed(0.00564971751412429377, 1, -nbits);
    elsif (x=178) then return to_sfixed(0.00561797752808988748, 1, -nbits);
    elsif (x=179) then return to_sfixed(0.00558659217877094990, 1, -nbits);
    elsif (x=180) then return to_sfixed(0.00555555555555555577, 1, -nbits);
    elsif (x=181) then return to_sfixed(0.00552486187845303844, 1, -nbits);
    elsif (x=182) then return to_sfixed(0.00549450549450549493, 1, -nbits);
    elsif (x=183) then return to_sfixed(0.00546448087431693989, 1, -nbits);
    elsif (x=184) then return to_sfixed(0.00543478260869565202, 1, -nbits);
    elsif (x=185) then return to_sfixed(0.00540540540540540571, 1, -nbits);
    elsif (x=186) then return to_sfixed(0.00537634408602150581, 1, -nbits);
    elsif (x=187) then return to_sfixed(0.00534759358288770022, 1, -nbits);
    elsif (x=188) then return to_sfixed(0.00531914893617021264, 1, -nbits);
    elsif (x=189) then return to_sfixed(0.00529100529100529071, 1, -nbits);
    elsif (x=190) then return to_sfixed(0.00526315789473684199, 1, -nbits);
    elsif (x=191) then return to_sfixed(0.00523560209424083801, 1, -nbits);
    elsif (x=192) then return to_sfixed(0.00520833333333333304, 1, -nbits);
    elsif (x=193) then return to_sfixed(0.00518134715025906755, 1, -nbits);
    elsif (x=194) then return to_sfixed(0.00515463917525773186, 1, -nbits);
    elsif (x=195) then return to_sfixed(0.00512820512820512820, 1, -nbits);
    elsif (x=196) then return to_sfixed(0.00510204081632653021, 1, -nbits);
    elsif (x=197) then return to_sfixed(0.00507614213197969504, 1, -nbits);
    elsif (x=198) then return to_sfixed(0.00505050505050505093, 1, -nbits);
    elsif (x=199) then return to_sfixed(0.00502512562814070359, 1, -nbits);
    elsif (x=200) then return to_sfixed(0.00500000000000000010, 1, -nbits);
    elsif (x=201) then return to_sfixed(0.00497512437810945264, 1, -nbits);
    elsif (x=202) then return to_sfixed(0.00495049504950495056, 1, -nbits);
    elsif (x=203) then return to_sfixed(0.00492610837438423651, 1, -nbits);
    elsif (x=204) then return to_sfixed(0.00490196078431372542, 1, -nbits);
    elsif (x=205) then return to_sfixed(0.00487804878048780487, 1, -nbits);
    elsif (x=206) then return to_sfixed(0.00485436893203883453, 1, -nbits);
    elsif (x=207) then return to_sfixed(0.00483091787439613504, 1, -nbits);
    elsif (x=208) then return to_sfixed(0.00480769230769230796, 1, -nbits);
    elsif (x=209) then return to_sfixed(0.00478468899521531082, 1, -nbits);
    elsif (x=210) then return to_sfixed(0.00476190476190476233, 1, -nbits);
    elsif (x=211) then return to_sfixed(0.00473933649289099562, 1, -nbits);
    elsif (x=212) then return to_sfixed(0.00471698113207547152, 1, -nbits);
    elsif (x=213) then return to_sfixed(0.00469483568075117381, 1, -nbits);
    elsif (x=214) then return to_sfixed(0.00467289719626168189, 1, -nbits);
    elsif (x=215) then return to_sfixed(0.00465116279069767435, 1, -nbits);
    elsif (x=216) then return to_sfixed(0.00462962962962962937, 1, -nbits);
    elsif (x=217) then return to_sfixed(0.00460829493087557603, 1, -nbits);
    elsif (x=218) then return to_sfixed(0.00458715596330275255, 1, -nbits);
    elsif (x=219) then return to_sfixed(0.00456621004566210020, 1, -nbits);
    elsif (x=220) then return to_sfixed(0.00454545454545454523, 1, -nbits);
    elsif (x=221) then return to_sfixed(0.00452488687782805470, 1, -nbits);
    elsif (x=222) then return to_sfixed(0.00450450450450450447, 1, -nbits);
    elsif (x=223) then return to_sfixed(0.00448430493273542594, 1, -nbits);
    elsif (x=224) then return to_sfixed(0.00446428571428571404, 1, -nbits);
    elsif (x=225) then return to_sfixed(0.00444444444444444444, 1, -nbits);
    elsif (x=226) then return to_sfixed(0.00442477876106194684, 1, -nbits);
    elsif (x=227) then return to_sfixed(0.00440528634361233521, 1, -nbits);
    elsif (x=228) then return to_sfixed(0.00438596491228070151, 1, -nbits);
    elsif (x=229) then return to_sfixed(0.00436681222707423558, 1, -nbits);
    elsif (x=230) then return to_sfixed(0.00434782608695652179, 1, -nbits);
    elsif (x=231) then return to_sfixed(0.00432900432900432900, 1, -nbits);
    elsif (x=232) then return to_sfixed(0.00431034482758620684, 1, -nbits);
    elsif (x=233) then return to_sfixed(0.00429184549356223174, 1, -nbits);
    elsif (x=234) then return to_sfixed(0.00427350427350427393, 1, -nbits);
    elsif (x=235) then return to_sfixed(0.00425531914893617028, 1, -nbits);
    elsif (x=236) then return to_sfixed(0.00423728813559322032, 1, -nbits);
    elsif (x=237) then return to_sfixed(0.00421940928270042159, 1, -nbits);
    elsif (x=238) then return to_sfixed(0.00420168067226890738, 1, -nbits);
    elsif (x=239) then return to_sfixed(0.00418410041841004148, 1, -nbits);
    elsif (x=240) then return to_sfixed(0.00416666666666666661, 1, -nbits);
    elsif (x=241) then return to_sfixed(0.00414937759336099585, 1, -nbits);
    elsif (x=242) then return to_sfixed(0.00413223140495867780, 1, -nbits);
    elsif (x=243) then return to_sfixed(0.00411522633744856002, 1, -nbits);
    elsif (x=244) then return to_sfixed(0.00409836065573770513, 1, -nbits);
    elsif (x=245) then return to_sfixed(0.00408163265306122486, 1, -nbits);
    elsif (x=246) then return to_sfixed(0.00406504065040650450, 1, -nbits);
    elsif (x=247) then return to_sfixed(0.00404858299595141705, 1, -nbits);
    elsif (x=248) then return to_sfixed(0.00403225806451612892, 1, -nbits);
    elsif (x=249) then return to_sfixed(0.00401606425702811208, 1, -nbits);
    elsif (x=250) then return to_sfixed(0.00400000000000000008, 1, -nbits);
    elsif (x=251) then return to_sfixed(0.00398406374501992025, 1, -nbits);
    elsif (x=252) then return to_sfixed(0.00396825396825396803, 1, -nbits);
    elsif (x=253) then return to_sfixed(0.00395256916996047404, 1, -nbits);
    elsif (x=254) then return to_sfixed(0.00393700787401574798, 1, -nbits);
    elsif (x=255) then return to_sfixed(0.00392156862745098034, 1, -nbits);
    elsif (x=256) then return to_sfixed(0.00390625000000000000, 1, -nbits);
    elsif (x=257) then return to_sfixed(0.00389105058365758760, 1, -nbits);
    elsif (x=258) then return to_sfixed(0.00387596899224806196, 1, -nbits);
    elsif (x=259) then return to_sfixed(0.00386100386100386109, 1, -nbits);
    elsif (x=260) then return to_sfixed(0.00384615384615384637, 1, -nbits);
    elsif (x=261) then return to_sfixed(0.00383141762452107260, 1, -nbits);
    elsif (x=262) then return to_sfixed(0.00381679389312977084, 1, -nbits);
    elsif (x=263) then return to_sfixed(0.00380228136882129275, 1, -nbits);
    elsif (x=264) then return to_sfixed(0.00378787878787878798, 1, -nbits);
    elsif (x=265) then return to_sfixed(0.00377358490566037739, 1, -nbits);
    elsif (x=266) then return to_sfixed(0.00375939849624060130, 1, -nbits);
    elsif (x=267) then return to_sfixed(0.00374531835205992513, 1, -nbits);
    elsif (x=268) then return to_sfixed(0.00373134328358208948, 1, -nbits);
    elsif (x=269) then return to_sfixed(0.00371747211895910763, 1, -nbits);
    elsif (x=270) then return to_sfixed(0.00370370370370370385, 1, -nbits);
    elsif (x=271) then return to_sfixed(0.00369003690036900358, 1, -nbits);
    elsif (x=272) then return to_sfixed(0.00367647058823529407, 1, -nbits);
    elsif (x=273) then return to_sfixed(0.00366300366300366300, 1, -nbits);
    elsif (x=274) then return to_sfixed(0.00364963503649635024, 1, -nbits);
    elsif (x=275) then return to_sfixed(0.00363636363636363636, 1, -nbits);
    elsif (x=276) then return to_sfixed(0.00362318840579710149, 1, -nbits);
    elsif (x=277) then return to_sfixed(0.00361010830324909760, 1, -nbits);
    elsif (x=278) then return to_sfixed(0.00359712230215827357, 1, -nbits);
    elsif (x=279) then return to_sfixed(0.00358422939068100358, 1, -nbits);
    elsif (x=280) then return to_sfixed(0.00357142857142857132, 1, -nbits);
    elsif (x=281) then return to_sfixed(0.00355871886120996423, 1, -nbits);
    elsif (x=282) then return to_sfixed(0.00354609929078014176, 1, -nbits);
    elsif (x=283) then return to_sfixed(0.00353356890459363953, 1, -nbits);
    elsif (x=284) then return to_sfixed(0.00352112676056338036, 1, -nbits);
    elsif (x=285) then return to_sfixed(0.00350877192982456147, 1, -nbits);
    elsif (x=286) then return to_sfixed(0.00349650349650349650, 1, -nbits);
    elsif (x=287) then return to_sfixed(0.00348432055749128920, 1, -nbits);
    elsif (x=288) then return to_sfixed(0.00347222222222222203, 1, -nbits);
    elsif (x=289) then return to_sfixed(0.00346020761245674751, 1, -nbits);
    elsif (x=290) then return to_sfixed(0.00344827586206896547, 1, -nbits);
    elsif (x=291) then return to_sfixed(0.00343642611683848791, 1, -nbits);
    elsif (x=292) then return to_sfixed(0.00342465753424657515, 1, -nbits);
    elsif (x=293) then return to_sfixed(0.00341296928327645055, 1, -nbits);
    elsif (x=294) then return to_sfixed(0.00340136054421768695, 1, -nbits);
    elsif (x=295) then return to_sfixed(0.00338983050847457617, 1, -nbits);
    elsif (x=296) then return to_sfixed(0.00337837837837837857, 1, -nbits);
    elsif (x=297) then return to_sfixed(0.00336700336700336686, 1, -nbits);
    elsif (x=298) then return to_sfixed(0.00335570469798657711, 1, -nbits);
    elsif (x=299) then return to_sfixed(0.00334448160535117051, 1, -nbits);
    elsif (x=300) then return to_sfixed(0.00333333333333333355, 1, -nbits);
    elsif (x=301) then return to_sfixed(0.00332225913621262466, 1, -nbits);
    elsif (x=302) then return to_sfixed(0.00331125827814569536, 1, -nbits);
    elsif (x=303) then return to_sfixed(0.00330033003300330037, 1, -nbits);
    elsif (x=304) then return to_sfixed(0.00328947368421052613, 1, -nbits);
    elsif (x=305) then return to_sfixed(0.00327868852459016393, 1, -nbits);
    elsif (x=306) then return to_sfixed(0.00326797385620915043, 1, -nbits);
    elsif (x=307) then return to_sfixed(0.00325732899022801317, 1, -nbits);
    elsif (x=308) then return to_sfixed(0.00324675324675324697, 1, -nbits);
    elsif (x=309) then return to_sfixed(0.00323624595469255679, 1, -nbits);
    elsif (x=310) then return to_sfixed(0.00322580645161290322, 1, -nbits);
    elsif (x=311) then return to_sfixed(0.00321543408360128614, 1, -nbits);
    elsif (x=312) then return to_sfixed(0.00320512820512820502, 1, -nbits);
    elsif (x=313) then return to_sfixed(0.00319488817891373789, 1, -nbits);
    elsif (x=314) then return to_sfixed(0.00318471337579617850, 1, -nbits);
    elsif (x=315) then return to_sfixed(0.00317460317460317460, 1, -nbits);
    elsif (x=316) then return to_sfixed(0.00316455696202531641, 1, -nbits);
    elsif (x=317) then return to_sfixed(0.00315457413249211347, 1, -nbits);
    elsif (x=318) then return to_sfixed(0.00314465408805031463, 1, -nbits);
    elsif (x=319) then return to_sfixed(0.00313479623824451398, 1, -nbits);
    elsif (x=320) then return to_sfixed(0.00312500000000000017, 1, -nbits);
    elsif (x=321) then return to_sfixed(0.00311526479750778807, 1, -nbits);
    elsif (x=322) then return to_sfixed(0.00310559006211180103, 1, -nbits);
    elsif (x=323) then return to_sfixed(0.00309597523219814260, 1, -nbits);
    elsif (x=324) then return to_sfixed(0.00308641975308641958, 1, -nbits);
    elsif (x=325) then return to_sfixed(0.00307692307692307692, 1, -nbits);
    elsif (x=326) then return to_sfixed(0.00306748466257668719, 1, -nbits);
    elsif (x=327) then return to_sfixed(0.00305810397553516822, 1, -nbits);
    elsif (x=328) then return to_sfixed(0.00304878048780487815, 1, -nbits);
    elsif (x=329) then return to_sfixed(0.00303951367781155014, 1, -nbits);
    elsif (x=330) then return to_sfixed(0.00303030303030303030, 1, -nbits);
    elsif (x=331) then return to_sfixed(0.00302114803625377643, 1, -nbits);
    elsif (x=332) then return to_sfixed(0.00301204819277108449, 1, -nbits);
    elsif (x=333) then return to_sfixed(0.00300300300300300298, 1, -nbits);
    elsif (x=334) then return to_sfixed(0.00299401197604790437, 1, -nbits);
    elsif (x=335) then return to_sfixed(0.00298507462686567167, 1, -nbits);
    elsif (x=336) then return to_sfixed(0.00297619047619047603, 1, -nbits);
    elsif (x=337) then return to_sfixed(0.00296735905044510397, 1, -nbits);
    elsif (x=338) then return to_sfixed(0.00295857988165680466, 1, -nbits);
    elsif (x=339) then return to_sfixed(0.00294985250737463123, 1, -nbits);
    elsif (x=340) then return to_sfixed(0.00294117647058823525, 1, -nbits);
    elsif (x=341) then return to_sfixed(0.00293255131964809384, 1, -nbits);
    elsif (x=342) then return to_sfixed(0.00292397660818713434, 1, -nbits);
    elsif (x=343) then return to_sfixed(0.00291545189504373173, 1, -nbits);
    elsif (x=344) then return to_sfixed(0.00290697674418604647, 1, -nbits);
    elsif (x=345) then return to_sfixed(0.00289855072463768119, 1, -nbits);
    elsif (x=346) then return to_sfixed(0.00289017341040462413, 1, -nbits);
    elsif (x=347) then return to_sfixed(0.00288184438040345802, 1, -nbits);
    elsif (x=348) then return to_sfixed(0.00287356321839080456, 1, -nbits);
    elsif (x=349) then return to_sfixed(0.00286532951289398272, 1, -nbits);
    elsif (x=350) then return to_sfixed(0.00285714285714285714, 1, -nbits);
    elsif (x=351) then return to_sfixed(0.00284900284900284914, 1, -nbits);
    elsif (x=352) then return to_sfixed(0.00284090909090909099, 1, -nbits);
    elsif (x=353) then return to_sfixed(0.00283286118980169985, 1, -nbits);
    elsif (x=354) then return to_sfixed(0.00282485875706214688, 1, -nbits);
    elsif (x=355) then return to_sfixed(0.00281690140845070438, 1, -nbits);
    elsif (x=356) then return to_sfixed(0.00280898876404494374, 1, -nbits);
    elsif (x=357) then return to_sfixed(0.00280112044817927173, 1, -nbits);
    elsif (x=358) then return to_sfixed(0.00279329608938547495, 1, -nbits);
    elsif (x=359) then return to_sfixed(0.00278551532033426185, 1, -nbits);
    elsif (x=360) then return to_sfixed(0.00277777777777777788, 1, -nbits);
    elsif (x=361) then return to_sfixed(0.00277008310249307480, 1, -nbits);
    elsif (x=362) then return to_sfixed(0.00276243093922651922, 1, -nbits);
    elsif (x=363) then return to_sfixed(0.00275482093663911853, 1, -nbits);
    elsif (x=364) then return to_sfixed(0.00274725274725274747, 1, -nbits);
    elsif (x=365) then return to_sfixed(0.00273972602739726030, 1, -nbits);
    elsif (x=366) then return to_sfixed(0.00273224043715846994, 1, -nbits);
    elsif (x=367) then return to_sfixed(0.00272479564032697538, 1, -nbits);
    elsif (x=368) then return to_sfixed(0.00271739130434782601, 1, -nbits);
    elsif (x=369) then return to_sfixed(0.00271002710027100271, 1, -nbits);
    elsif (x=370) then return to_sfixed(0.00270270270270270285, 1, -nbits);
    elsif (x=371) then return to_sfixed(0.00269541778975741254, 1, -nbits);
    elsif (x=372) then return to_sfixed(0.00268817204301075290, 1, -nbits);
    elsif (x=373) then return to_sfixed(0.00268096514745308316, 1, -nbits);
    elsif (x=374) then return to_sfixed(0.00267379679144385011, 1, -nbits);
    elsif (x=375) then return to_sfixed(0.00266666666666666658, 1, -nbits);
    elsif (x=376) then return to_sfixed(0.00265957446808510632, 1, -nbits);
    elsif (x=377) then return to_sfixed(0.00265251989389920411, 1, -nbits);
    elsif (x=378) then return to_sfixed(0.00264550264550264536, 1, -nbits);
    elsif (x=379) then return to_sfixed(0.00263852242744063315, 1, -nbits);
    elsif (x=380) then return to_sfixed(0.00263157894736842099, 1, -nbits);
    elsif (x=381) then return to_sfixed(0.00262467191601049865, 1, -nbits);
    elsif (x=382) then return to_sfixed(0.00261780104712041901, 1, -nbits);
    elsif (x=383) then return to_sfixed(0.00261096605744125330, 1, -nbits);
    elsif (x=384) then return to_sfixed(0.00260416666666666652, 1, -nbits);
    elsif (x=385) then return to_sfixed(0.00259740259740259740, 1, -nbits);
    elsif (x=386) then return to_sfixed(0.00259067357512953378, 1, -nbits);
    elsif (x=387) then return to_sfixed(0.00258397932816537479, 1, -nbits);
    elsif (x=388) then return to_sfixed(0.00257731958762886593, 1, -nbits);
    elsif (x=389) then return to_sfixed(0.00257069408740359879, 1, -nbits);
    elsif (x=390) then return to_sfixed(0.00256410256410256410, 1, -nbits);
    elsif (x=391) then return to_sfixed(0.00255754475703324829, 1, -nbits);
    elsif (x=392) then return to_sfixed(0.00255102040816326510, 1, -nbits);
    elsif (x=393) then return to_sfixed(0.00254452926208651418, 1, -nbits);
    elsif (x=394) then return to_sfixed(0.00253807106598984752, 1, -nbits);
    elsif (x=395) then return to_sfixed(0.00253164556962025321, 1, -nbits);
    elsif (x=396) then return to_sfixed(0.00252525252525252547, 1, -nbits);
    elsif (x=397) then return to_sfixed(0.00251889168765743066, 1, -nbits);
    elsif (x=398) then return to_sfixed(0.00251256281407035180, 1, -nbits);
    elsif (x=399) then return to_sfixed(0.00250626566416040086, 1, -nbits);
    elsif (x=400) then return to_sfixed(0.00250000000000000005, 1, -nbits);
    elsif (x=401) then return to_sfixed(0.00249376558603491266, 1, -nbits);
    elsif (x=402) then return to_sfixed(0.00248756218905472632, 1, -nbits);
    elsif (x=403) then return to_sfixed(0.00248138957816377171, 1, -nbits);
    elsif (x=404) then return to_sfixed(0.00247524752475247528, 1, -nbits);
    elsif (x=405) then return to_sfixed(0.00246913580246913575, 1, -nbits);
    elsif (x=406) then return to_sfixed(0.00246305418719211825, 1, -nbits);
    elsif (x=407) then return to_sfixed(0.00245700245700245694, 1, -nbits);
    elsif (x=408) then return to_sfixed(0.00245098039215686271, 1, -nbits);
    elsif (x=409) then return to_sfixed(0.00244498777506112468, 1, -nbits);
    elsif (x=410) then return to_sfixed(0.00243902439024390244, 1, -nbits);
    elsif (x=411) then return to_sfixed(0.00243309002433090031, 1, -nbits);
    elsif (x=412) then return to_sfixed(0.00242718446601941727, 1, -nbits);
    elsif (x=413) then return to_sfixed(0.00242130750605326888, 1, -nbits);
    elsif (x=414) then return to_sfixed(0.00241545893719806752, 1, -nbits);
    elsif (x=415) then return to_sfixed(0.00240963855421686768, 1, -nbits);
    elsif (x=416) then return to_sfixed(0.00240384615384615398, 1, -nbits);
    elsif (x=417) then return to_sfixed(0.00239808153477218209, 1, -nbits);
    elsif (x=418) then return to_sfixed(0.00239234449760765541, 1, -nbits);
    elsif (x=419) then return to_sfixed(0.00238663484486873519, 1, -nbits);
    elsif (x=420) then return to_sfixed(0.00238095238095238117, 1, -nbits);
    elsif (x=421) then return to_sfixed(0.00237529691211401436, 1, -nbits);
    elsif (x=422) then return to_sfixed(0.00236966824644549781, 1, -nbits);
    elsif (x=423) then return to_sfixed(0.00236406619385342784, 1, -nbits);
    elsif (x=424) then return to_sfixed(0.00235849056603773576, 1, -nbits);
    elsif (x=425) then return to_sfixed(0.00235294117647058803, 1, -nbits);
    elsif (x=426) then return to_sfixed(0.00234741784037558691, 1, -nbits);
    elsif (x=427) then return to_sfixed(0.00234192037470725995, 1, -nbits);
    elsif (x=428) then return to_sfixed(0.00233644859813084095, 1, -nbits);
    elsif (x=429) then return to_sfixed(0.00233100233100233100, 1, -nbits);
    elsif (x=430) then return to_sfixed(0.00232558139534883718, 1, -nbits);
    elsif (x=431) then return to_sfixed(0.00232018561484918784, 1, -nbits);
    elsif (x=432) then return to_sfixed(0.00231481481481481469, 1, -nbits);
    elsif (x=433) then return to_sfixed(0.00230946882217090066, 1, -nbits);
    elsif (x=434) then return to_sfixed(0.00230414746543778802, 1, -nbits);
    elsif (x=435) then return to_sfixed(0.00229885057471264365, 1, -nbits);
    elsif (x=436) then return to_sfixed(0.00229357798165137627, 1, -nbits);
    elsif (x=437) then return to_sfixed(0.00228832951945080092, 1, -nbits);
    elsif (x=438) then return to_sfixed(0.00228310502283105010, 1, -nbits);
    elsif (x=439) then return to_sfixed(0.00227790432801822313, 1, -nbits);
    elsif (x=440) then return to_sfixed(0.00227272727272727262, 1, -nbits);
    elsif (x=441) then return to_sfixed(0.00226757369614512478, 1, -nbits);
    elsif (x=442) then return to_sfixed(0.00226244343891402735, 1, -nbits);
    elsif (x=443) then return to_sfixed(0.00225733634311512396, 1, -nbits);
    elsif (x=444) then return to_sfixed(0.00225225225225225223, 1, -nbits);
    elsif (x=445) then return to_sfixed(0.00224719101123595525, 1, -nbits);
    elsif (x=446) then return to_sfixed(0.00224215246636771297, 1, -nbits);
    elsif (x=447) then return to_sfixed(0.00223713646532438474, 1, -nbits);
    elsif (x=448) then return to_sfixed(0.00223214285714285702, 1, -nbits);
    elsif (x=449) then return to_sfixed(0.00222717149220489968, 1, -nbits);
    elsif (x=450) then return to_sfixed(0.00222222222222222222, 1, -nbits);
    elsif (x=451) then return to_sfixed(0.00221729490022172949, 1, -nbits);
    elsif (x=452) then return to_sfixed(0.00221238938053097342, 1, -nbits);
    elsif (x=453) then return to_sfixed(0.00220750551876379691, 1, -nbits);
    elsif (x=454) then return to_sfixed(0.00220264317180616761, 1, -nbits);
    elsif (x=455) then return to_sfixed(0.00219780219780219780, 1, -nbits);
    elsif (x=456) then return to_sfixed(0.00219298245614035076, 1, -nbits);
    elsif (x=457) then return to_sfixed(0.00218818380743982487, 1, -nbits);
    elsif (x=458) then return to_sfixed(0.00218340611353711779, 1, -nbits);
    elsif (x=459) then return to_sfixed(0.00217864923747276710, 1, -nbits);
    elsif (x=460) then return to_sfixed(0.00217391304347826090, 1, -nbits);
    elsif (x=461) then return to_sfixed(0.00216919739696312371, 1, -nbits);
    elsif (x=462) then return to_sfixed(0.00216450216450216450, 1, -nbits);
    elsif (x=463) then return to_sfixed(0.00215982721382289430, 1, -nbits);
    elsif (x=464) then return to_sfixed(0.00215517241379310342, 1, -nbits);
    elsif (x=465) then return to_sfixed(0.00215053763440860215, 1, -nbits);
    elsif (x=466) then return to_sfixed(0.00214592274678111587, 1, -nbits);
    elsif (x=467) then return to_sfixed(0.00214132762312633845, 1, -nbits);
    elsif (x=468) then return to_sfixed(0.00213675213675213697, 1, -nbits);
    elsif (x=469) then return to_sfixed(0.00213219616204690827, 1, -nbits);
    elsif (x=470) then return to_sfixed(0.00212765957446808514, 1, -nbits);
    elsif (x=471) then return to_sfixed(0.00212314225053078552, 1, -nbits);
    elsif (x=472) then return to_sfixed(0.00211864406779661016, 1, -nbits);
    elsif (x=473) then return to_sfixed(0.00211416490486257937, 1, -nbits);
    elsif (x=474) then return to_sfixed(0.00210970464135021079, 1, -nbits);
    elsif (x=475) then return to_sfixed(0.00210526315789473679, 1, -nbits);
    elsif (x=476) then return to_sfixed(0.00210084033613445369, 1, -nbits);
    elsif (x=477) then return to_sfixed(0.00209643605870020976, 1, -nbits);
    elsif (x=478) then return to_sfixed(0.00209205020920502074, 1, -nbits);
    elsif (x=479) then return to_sfixed(0.00208768267223382025, 1, -nbits);
    elsif (x=480) then return to_sfixed(0.00208333333333333330, 1, -nbits);
    elsif (x=481) then return to_sfixed(0.00207900207900207912, 1, -nbits);
    elsif (x=482) then return to_sfixed(0.00207468879668049793, 1, -nbits);
    elsif (x=483) then return to_sfixed(0.00207039337474120098, 1, -nbits);
    elsif (x=484) then return to_sfixed(0.00206611570247933890, 1, -nbits);
    elsif (x=485) then return to_sfixed(0.00206185567010309283, 1, -nbits);
    elsif (x=486) then return to_sfixed(0.00205761316872428001, 1, -nbits);
    elsif (x=487) then return to_sfixed(0.00205338809034907605, 1, -nbits);
    elsif (x=488) then return to_sfixed(0.00204918032786885257, 1, -nbits);
    elsif (x=489) then return to_sfixed(0.00204498977505112494, 1, -nbits);
    elsif (x=490) then return to_sfixed(0.00204081632653061243, 1, -nbits);
    elsif (x=491) then return to_sfixed(0.00203665987780040714, 1, -nbits);
    elsif (x=492) then return to_sfixed(0.00203252032520325225, 1, -nbits);
    elsif (x=493) then return to_sfixed(0.00202839756592292086, 1, -nbits);
    elsif (x=494) then return to_sfixed(0.00202429149797570852, 1, -nbits);
    elsif (x=495) then return to_sfixed(0.00202020202020202020, 1, -nbits);
    elsif (x=496) then return to_sfixed(0.00201612903225806446, 1, -nbits);
    elsif (x=497) then return to_sfixed(0.00201207243460764604, 1, -nbits);
    elsif (x=498) then return to_sfixed(0.00200803212851405604, 1, -nbits);
    elsif (x=499) then return to_sfixed(0.00200400801603206396, 1, -nbits);
    elsif (x=500) then return to_sfixed(0.00200000000000000004, 1, -nbits);
    elsif (x=501) then return to_sfixed(0.00199600798403193596, 1, -nbits);
    elsif (x=502) then return to_sfixed(0.00199203187250996012, 1, -nbits);
    elsif (x=503) then return to_sfixed(0.00198807157057654055, 1, -nbits);
    elsif (x=504) then return to_sfixed(0.00198412698412698402, 1, -nbits);
    elsif (x=505) then return to_sfixed(0.00198019801980198022, 1, -nbits);
    elsif (x=506) then return to_sfixed(0.00197628458498023702, 1, -nbits);
    elsif (x=507) then return to_sfixed(0.00197238658777120325, 1, -nbits);
    elsif (x=508) then return to_sfixed(0.00196850393700787399, 1, -nbits);
    elsif (x=509) then return to_sfixed(0.00196463654223968552, 1, -nbits);
    elsif (x=510) then return to_sfixed(0.00196078431372549017, 1, -nbits);
    elsif (x=511) then return to_sfixed(0.00195694716242661437, 1, -nbits);
    elsif (x=512) then return to_sfixed(0.00195312500000000000, 1, -nbits);
    elsif (x=513) then return to_sfixed(0.00194931773879142289, 1, -nbits);
    elsif (x=514) then return to_sfixed(0.00194552529182879380, 1, -nbits);
    elsif (x=515) then return to_sfixed(0.00194174757281553390, 1, -nbits);
    elsif (x=516) then return to_sfixed(0.00193798449612403098, 1, -nbits);
    elsif (x=517) then return to_sfixed(0.00193423597678916829, 1, -nbits);
    elsif (x=518) then return to_sfixed(0.00193050193050193055, 1, -nbits);
    elsif (x=519) then return to_sfixed(0.00192678227360308283, 1, -nbits);
    elsif (x=520) then return to_sfixed(0.00192307692307692318, 1, -nbits);
    elsif (x=521) then return to_sfixed(0.00191938579654510550, 1, -nbits);
    elsif (x=522) then return to_sfixed(0.00191570881226053630, 1, -nbits);
    elsif (x=523) then return to_sfixed(0.00191204588910133836, 1, -nbits);
    elsif (x=524) then return to_sfixed(0.00190839694656488542, 1, -nbits);
    elsif (x=525) then return to_sfixed(0.00190476190476190476, 1, -nbits);
    elsif (x=526) then return to_sfixed(0.00190114068441064638, 1, -nbits);
    elsif (x=527) then return to_sfixed(0.00189753320683111958, 1, -nbits);
    elsif (x=528) then return to_sfixed(0.00189393939393939399, 1, -nbits);
    elsif (x=529) then return to_sfixed(0.00189035916824196602, 1, -nbits);
    elsif (x=530) then return to_sfixed(0.00188679245283018869, 1, -nbits);
    elsif (x=531) then return to_sfixed(0.00188323917137476452, 1, -nbits);
    elsif (x=532) then return to_sfixed(0.00187969924812030065, 1, -nbits);
    elsif (x=533) then return to_sfixed(0.00187617260787992495, 1, -nbits);
    elsif (x=534) then return to_sfixed(0.00187265917602996257, 1, -nbits);
    elsif (x=535) then return to_sfixed(0.00186915887850467297, 1, -nbits);
    elsif (x=536) then return to_sfixed(0.00186567164179104474, 1, -nbits);
    elsif (x=537) then return to_sfixed(0.00186219739292364989, 1, -nbits);
    elsif (x=538) then return to_sfixed(0.00185873605947955382, 1, -nbits);
    elsif (x=539) then return to_sfixed(0.00185528756957328389, 1, -nbits);
    elsif (x=540) then return to_sfixed(0.00185185185185185192, 1, -nbits);
    elsif (x=541) then return to_sfixed(0.00184842883548983362, 1, -nbits);
    elsif (x=542) then return to_sfixed(0.00184501845018450179, 1, -nbits);
    elsif (x=543) then return to_sfixed(0.00184162062615101296, 1, -nbits);
    elsif (x=544) then return to_sfixed(0.00183823529411764703, 1, -nbits);
    elsif (x=545) then return to_sfixed(0.00183486238532110102, 1, -nbits);
    elsif (x=546) then return to_sfixed(0.00183150183150183150, 1, -nbits);
    elsif (x=547) then return to_sfixed(0.00182815356489945155, 1, -nbits);
    elsif (x=548) then return to_sfixed(0.00182481751824817512, 1, -nbits);
    elsif (x=549) then return to_sfixed(0.00182149362477231330, 1, -nbits);
    elsif (x=550) then return to_sfixed(0.00181818181818181818, 1, -nbits);
    elsif (x=551) then return to_sfixed(0.00181488203266787652, 1, -nbits);
    elsif (x=552) then return to_sfixed(0.00181159420289855075, 1, -nbits);
    elsif (x=553) then return to_sfixed(0.00180831826401446649, 1, -nbits);
    elsif (x=554) then return to_sfixed(0.00180505415162454880, 1, -nbits);
    elsif (x=555) then return to_sfixed(0.00180180180180180183, 1, -nbits);
    elsif (x=556) then return to_sfixed(0.00179856115107913678, 1, -nbits);
    elsif (x=557) then return to_sfixed(0.00179533213644524244, 1, -nbits);
    elsif (x=558) then return to_sfixed(0.00179211469534050179, 1, -nbits);
    elsif (x=559) then return to_sfixed(0.00178890876565295171, 1, -nbits);
    elsif (x=560) then return to_sfixed(0.00178571428571428566, 1, -nbits);
    elsif (x=561) then return to_sfixed(0.00178253119429590007, 1, -nbits);
    elsif (x=562) then return to_sfixed(0.00177935943060498212, 1, -nbits);
    elsif (x=563) then return to_sfixed(0.00177619893428063950, 1, -nbits);
    elsif (x=564) then return to_sfixed(0.00177304964539007088, 1, -nbits);
    elsif (x=565) then return to_sfixed(0.00176991150442477874, 1, -nbits);
    elsif (x=566) then return to_sfixed(0.00176678445229681976, 1, -nbits);
    elsif (x=567) then return to_sfixed(0.00176366843033509690, 1, -nbits);
    elsif (x=568) then return to_sfixed(0.00176056338028169018, 1, -nbits);
    elsif (x=569) then return to_sfixed(0.00175746924428822485, 1, -nbits);
    elsif (x=570) then return to_sfixed(0.00175438596491228073, 1, -nbits);
    elsif (x=571) then return to_sfixed(0.00175131348511383539, 1, -nbits);
    elsif (x=572) then return to_sfixed(0.00174825174825174825, 1, -nbits);
    elsif (x=573) then return to_sfixed(0.00174520069808027927, 1, -nbits);
    elsif (x=574) then return to_sfixed(0.00174216027874564460, 1, -nbits);
    elsif (x=575) then return to_sfixed(0.00173913043478260876, 1, -nbits);
    elsif (x=576) then return to_sfixed(0.00173611111111111101, 1, -nbits);
    elsif (x=577) then return to_sfixed(0.00173310225303292885, 1, -nbits);
    elsif (x=578) then return to_sfixed(0.00173010380622837375, 1, -nbits);
    elsif (x=579) then return to_sfixed(0.00172711571675302237, 1, -nbits);
    elsif (x=580) then return to_sfixed(0.00172413793103448273, 1, -nbits);
    elsif (x=581) then return to_sfixed(0.00172117039586919111, 1, -nbits);
    elsif (x=582) then return to_sfixed(0.00171821305841924395, 1, -nbits);
    elsif (x=583) then return to_sfixed(0.00171526586620926241, 1, -nbits);
    elsif (x=584) then return to_sfixed(0.00171232876712328758, 1, -nbits);
    elsif (x=585) then return to_sfixed(0.00170940170940170940, 1, -nbits);
    elsif (x=586) then return to_sfixed(0.00170648464163822527, 1, -nbits);
    elsif (x=587) then return to_sfixed(0.00170357751277683137, 1, -nbits);
    elsif (x=588) then return to_sfixed(0.00170068027210884347, 1, -nbits);
    elsif (x=589) then return to_sfixed(0.00169779286926994904, 1, -nbits);
    elsif (x=590) then return to_sfixed(0.00169491525423728809, 1, -nbits);
    elsif (x=591) then return to_sfixed(0.00169204737732656508, 1, -nbits);
    elsif (x=592) then return to_sfixed(0.00168918918918918928, 1, -nbits);
    elsif (x=593) then return to_sfixed(0.00168634064080944342, 1, -nbits);
    elsif (x=594) then return to_sfixed(0.00168350168350168343, 1, -nbits);
    elsif (x=595) then return to_sfixed(0.00168067226890756313, 1, -nbits);
    elsif (x=596) then return to_sfixed(0.00167785234899328855, 1, -nbits);
    elsif (x=597) then return to_sfixed(0.00167504187604690120, 1, -nbits);
    elsif (x=598) then return to_sfixed(0.00167224080267558525, 1, -nbits);
    elsif (x=599) then return to_sfixed(0.00166944908180300506, 1, -nbits);
    elsif (x=600) then return to_sfixed(0.00166666666666666677, 1, -nbits);
    elsif (x=601) then return to_sfixed(0.00166389351081530786, 1, -nbits);
    elsif (x=602) then return to_sfixed(0.00166112956810631233, 1, -nbits);
    elsif (x=603) then return to_sfixed(0.00165837479270315095, 1, -nbits);
    elsif (x=604) then return to_sfixed(0.00165562913907284768, 1, -nbits);
    elsif (x=605) then return to_sfixed(0.00165289256198347103, 1, -nbits);
    elsif (x=606) then return to_sfixed(0.00165016501650165019, 1, -nbits);
    elsif (x=607) then return to_sfixed(0.00164744645799011534, 1, -nbits);
    elsif (x=608) then return to_sfixed(0.00164473684210526307, 1, -nbits);
    elsif (x=609) then return to_sfixed(0.00164203612479474543, 1, -nbits);
    elsif (x=610) then return to_sfixed(0.00163934426229508197, 1, -nbits);
    elsif (x=611) then return to_sfixed(0.00163666121112929631, 1, -nbits);
    elsif (x=612) then return to_sfixed(0.00163398692810457521, 1, -nbits);
    elsif (x=613) then return to_sfixed(0.00163132137030995114, 1, -nbits);
    elsif (x=614) then return to_sfixed(0.00162866449511400659, 1, -nbits);
    elsif (x=615) then return to_sfixed(0.00162601626016260162, 1, -nbits);
    elsif (x=616) then return to_sfixed(0.00162337662337662348, 1, -nbits);
    elsif (x=617) then return to_sfixed(0.00162074554294975681, 1, -nbits);
    elsif (x=618) then return to_sfixed(0.00161812297734627839, 1, -nbits);
    elsif (x=619) then return to_sfixed(0.00161550888529886924, 1, -nbits);
    elsif (x=620) then return to_sfixed(0.00161290322580645161, 1, -nbits);
    elsif (x=621) then return to_sfixed(0.00161030595813204508, 1, -nbits);
    elsif (x=622) then return to_sfixed(0.00160771704180064307, 1, -nbits);
    elsif (x=623) then return to_sfixed(0.00160513643659711074, 1, -nbits);
    elsif (x=624) then return to_sfixed(0.00160256410256410251, 1, -nbits);
    elsif (x=625) then return to_sfixed(0.00160000000000000008, 1, -nbits);
    elsif (x=626) then return to_sfixed(0.00159744408945686894, 1, -nbits);
    elsif (x=627) then return to_sfixed(0.00159489633173843701, 1, -nbits);
    elsif (x=628) then return to_sfixed(0.00159235668789808925, 1, -nbits);
    elsif (x=629) then return to_sfixed(0.00158982511923688404, 1, -nbits);
    elsif (x=630) then return to_sfixed(0.00158730158730158730, 1, -nbits);
    elsif (x=631) then return to_sfixed(0.00158478605388272589, 1, -nbits);
    elsif (x=632) then return to_sfixed(0.00158227848101265820, 1, -nbits);
    elsif (x=633) then return to_sfixed(0.00157977883096366506, 1, -nbits);
    elsif (x=634) then return to_sfixed(0.00157728706624605673, 1, -nbits);
    elsif (x=635) then return to_sfixed(0.00157480314960629919, 1, -nbits);
    elsif (x=636) then return to_sfixed(0.00157232704402515732, 1, -nbits);
    elsif (x=637) then return to_sfixed(0.00156985871271585566, 1, -nbits);
    elsif (x=638) then return to_sfixed(0.00156739811912225699, 1, -nbits);
    elsif (x=639) then return to_sfixed(0.00156494522691705794, 1, -nbits);
    elsif (x=640) then return to_sfixed(0.00156250000000000009, 1, -nbits);
    elsif (x=641) then return to_sfixed(0.00156006240249609990, 1, -nbits);
    elsif (x=642) then return to_sfixed(0.00155763239875389404, 1, -nbits);
    elsif (x=643) then return to_sfixed(0.00155520995334370140, 1, -nbits);
    elsif (x=644) then return to_sfixed(0.00155279503105590052, 1, -nbits);
    elsif (x=645) then return to_sfixed(0.00155038759689922478, 1, -nbits);
    elsif (x=646) then return to_sfixed(0.00154798761609907130, 1, -nbits);
    elsif (x=647) then return to_sfixed(0.00154559505409582686, 1, -nbits);
    elsif (x=648) then return to_sfixed(0.00154320987654320979, 1, -nbits);
    elsif (x=649) then return to_sfixed(0.00154083204930662563, 1, -nbits);
    elsif (x=650) then return to_sfixed(0.00153846153846153846, 1, -nbits);
    elsif (x=651) then return to_sfixed(0.00153609831029185868, 1, -nbits);
    elsif (x=652) then return to_sfixed(0.00153374233128834359, 1, -nbits);
    elsif (x=653) then return to_sfixed(0.00153139356814701384, 1, -nbits);
    elsif (x=654) then return to_sfixed(0.00152905198776758411, 1, -nbits);
    elsif (x=655) then return to_sfixed(0.00152671755725190838, 1, -nbits);
    elsif (x=656) then return to_sfixed(0.00152439024390243908, 1, -nbits);
    elsif (x=657) then return to_sfixed(0.00152207001522070007, 1, -nbits);
    elsif (x=658) then return to_sfixed(0.00151975683890577507, 1, -nbits);
    elsif (x=659) then return to_sfixed(0.00151745068285280733, 1, -nbits);
    elsif (x=660) then return to_sfixed(0.00151515151515151515, 1, -nbits);
    elsif (x=661) then return to_sfixed(0.00151285930408472016, 1, -nbits);
    elsif (x=662) then return to_sfixed(0.00151057401812688822, 1, -nbits);
    elsif (x=663) then return to_sfixed(0.00150829562594268483, 1, -nbits);
    elsif (x=664) then return to_sfixed(0.00150602409638554225, 1, -nbits);
    elsif (x=665) then return to_sfixed(0.00150375939849624069, 1, -nbits);
    elsif (x=666) then return to_sfixed(0.00150150150150150149, 1, -nbits);
    elsif (x=667) then return to_sfixed(0.00149925037481259365, 1, -nbits);
    elsif (x=668) then return to_sfixed(0.00149700598802395219, 1, -nbits);
    elsif (x=669) then return to_sfixed(0.00149476831091180872, 1, -nbits);
    elsif (x=670) then return to_sfixed(0.00149253731343283584, 1, -nbits);
    elsif (x=671) then return to_sfixed(0.00149031296572280179, 1, -nbits);
    elsif (x=672) then return to_sfixed(0.00148809523809523801, 1, -nbits);
    elsif (x=673) then return to_sfixed(0.00148588410104011880, 1, -nbits);
    elsif (x=674) then return to_sfixed(0.00148367952522255198, 1, -nbits);
    elsif (x=675) then return to_sfixed(0.00148148148148148141, 1, -nbits);
    elsif (x=676) then return to_sfixed(0.00147928994082840233, 1, -nbits);
    elsif (x=677) then return to_sfixed(0.00147710487444608577, 1, -nbits);
    elsif (x=678) then return to_sfixed(0.00147492625368731561, 1, -nbits);
    elsif (x=679) then return to_sfixed(0.00147275405007363767, 1, -nbits);
    elsif (x=680) then return to_sfixed(0.00147058823529411763, 1, -nbits);
    elsif (x=681) then return to_sfixed(0.00146842878120411152, 1, -nbits);
    elsif (x=682) then return to_sfixed(0.00146627565982404692, 1, -nbits);
    elsif (x=683) then return to_sfixed(0.00146412884333821380, 1, -nbits);
    elsif (x=684) then return to_sfixed(0.00146198830409356717, 1, -nbits);
    elsif (x=685) then return to_sfixed(0.00145985401459854005, 1, -nbits);
    elsif (x=686) then return to_sfixed(0.00145772594752186587, 1, -nbits);
    elsif (x=687) then return to_sfixed(0.00145560407569141200, 1, -nbits);
    elsif (x=688) then return to_sfixed(0.00145348837209302324, 1, -nbits);
    elsif (x=689) then return to_sfixed(0.00145137880986937590, 1, -nbits);
    elsif (x=690) then return to_sfixed(0.00144927536231884060, 1, -nbits);
    elsif (x=691) then return to_sfixed(0.00144717800289435590, 1, -nbits);
    elsif (x=692) then return to_sfixed(0.00144508670520231207, 1, -nbits);
    elsif (x=693) then return to_sfixed(0.00144300144300144300, 1, -nbits);
    elsif (x=694) then return to_sfixed(0.00144092219020172901, 1, -nbits);
    elsif (x=695) then return to_sfixed(0.00143884892086330938, 1, -nbits);
    elsif (x=696) then return to_sfixed(0.00143678160919540228, 1, -nbits);
    elsif (x=697) then return to_sfixed(0.00143472022955523680, 1, -nbits);
    elsif (x=698) then return to_sfixed(0.00143266475644699136, 1, -nbits);
    elsif (x=699) then return to_sfixed(0.00143061516452074391, 1, -nbits);
    elsif (x=700) then return to_sfixed(0.00142857142857142857, 1, -nbits);
    elsif (x=701) then return to_sfixed(0.00142653352353780318, 1, -nbits);
    elsif (x=702) then return to_sfixed(0.00142450142450142457, 1, -nbits);
    elsif (x=703) then return to_sfixed(0.00142247510668563307, 1, -nbits);
    elsif (x=704) then return to_sfixed(0.00142045454545454549, 1, -nbits);
    elsif (x=705) then return to_sfixed(0.00141843971631205683, 1, -nbits);
    elsif (x=706) then return to_sfixed(0.00141643059490084993, 1, -nbits);
    elsif (x=707) then return to_sfixed(0.00141442715700141448, 1, -nbits);
    elsif (x=708) then return to_sfixed(0.00141242937853107344, 1, -nbits);
    elsif (x=709) then return to_sfixed(0.00141043723554301831, 1, -nbits);
    elsif (x=710) then return to_sfixed(0.00140845070422535219, 1, -nbits);
    elsif (x=711) then return to_sfixed(0.00140646976090014067, 1, -nbits);
    elsif (x=712) then return to_sfixed(0.00140449438202247187, 1, -nbits);
    elsif (x=713) then return to_sfixed(0.00140252454417952310, 1, -nbits);
    elsif (x=714) then return to_sfixed(0.00140056022408963587, 1, -nbits);
    elsif (x=715) then return to_sfixed(0.00139860139860139860, 1, -nbits);
    elsif (x=716) then return to_sfixed(0.00139664804469273747, 1, -nbits);
    elsif (x=717) then return to_sfixed(0.00139470013947001390, 1, -nbits);
    elsif (x=718) then return to_sfixed(0.00139275766016713092, 1, -nbits);
    elsif (x=719) then return to_sfixed(0.00139082058414464528, 1, -nbits);
    elsif (x=720) then return to_sfixed(0.00138888888888888894, 1, -nbits);
    elsif (x=721) then return to_sfixed(0.00138696255201109574, 1, -nbits);
    elsif (x=722) then return to_sfixed(0.00138504155124653740, 1, -nbits);
    elsif (x=723) then return to_sfixed(0.00138312586445366536, 1, -nbits);
    elsif (x=724) then return to_sfixed(0.00138121546961325961, 1, -nbits);
    elsif (x=725) then return to_sfixed(0.00137931034482758610, 1, -nbits);
    elsif (x=726) then return to_sfixed(0.00137741046831955927, 1, -nbits);
    elsif (x=727) then return to_sfixed(0.00137551581843191198, 1, -nbits);
    elsif (x=728) then return to_sfixed(0.00137362637362637373, 1, -nbits);
    elsif (x=729) then return to_sfixed(0.00137174211248285312, 1, -nbits);
    elsif (x=730) then return to_sfixed(0.00136986301369863015, 1, -nbits);
    elsif (x=731) then return to_sfixed(0.00136798905608755128, 1, -nbits);
    elsif (x=732) then return to_sfixed(0.00136612021857923497, 1, -nbits);
    elsif (x=733) then return to_sfixed(0.00136425648021828104, 1, -nbits);
    elsif (x=734) then return to_sfixed(0.00136239782016348769, 1, -nbits);
    elsif (x=735) then return to_sfixed(0.00136054421768707474, 1, -nbits);
    elsif (x=736) then return to_sfixed(0.00135869565217391301, 1, -nbits);
    elsif (x=737) then return to_sfixed(0.00135685210312075973, 1, -nbits);
    elsif (x=738) then return to_sfixed(0.00135501355013550135, 1, -nbits);
    elsif (x=739) then return to_sfixed(0.00135317997293640064, 1, -nbits);
    elsif (x=740) then return to_sfixed(0.00135135135135135143, 1, -nbits);
    elsif (x=741) then return to_sfixed(0.00134952766531713894, 1, -nbits);
    elsif (x=742) then return to_sfixed(0.00134770889487870627, 1, -nbits);
    elsif (x=743) then return to_sfixed(0.00134589502018842531, 1, -nbits);
    elsif (x=744) then return to_sfixed(0.00134408602150537645, 1, -nbits);
    elsif (x=745) then return to_sfixed(0.00134228187919463080, 1, -nbits);
    elsif (x=746) then return to_sfixed(0.00134048257372654158, 1, -nbits);
    elsif (x=747) then return to_sfixed(0.00133868808567603743, 1, -nbits);
    elsif (x=748) then return to_sfixed(0.00133689839572192506, 1, -nbits);
    elsif (x=749) then return to_sfixed(0.00133511348464619489, 1, -nbits);
    elsif (x=750) then return to_sfixed(0.00133333333333333329, 1, -nbits);
    elsif (x=751) then return to_sfixed(0.00133155792276964057, 1, -nbits);
    elsif (x=752) then return to_sfixed(0.00132978723404255316, 1, -nbits);
    elsif (x=753) then return to_sfixed(0.00132802124833997334, 1, -nbits);
    elsif (x=754) then return to_sfixed(0.00132625994694960205, 1, -nbits);
    elsif (x=755) then return to_sfixed(0.00132450331125827814, 1, -nbits);
    elsif (x=756) then return to_sfixed(0.00132275132275132268, 1, -nbits);
    elsif (x=757) then return to_sfixed(0.00132100396301188905, 1, -nbits);
    elsif (x=758) then return to_sfixed(0.00131926121372031658, 1, -nbits);
    elsif (x=759) then return to_sfixed(0.00131752305665349149, 1, -nbits);
    elsif (x=760) then return to_sfixed(0.00131578947368421050, 1, -nbits);
    elsif (x=761) then return to_sfixed(0.00131406044678055193, 1, -nbits);
    elsif (x=762) then return to_sfixed(0.00131233595800524933, 1, -nbits);
    elsif (x=763) then return to_sfixed(0.00131061598951507209, 1, -nbits);
    elsif (x=764) then return to_sfixed(0.00130890052356020950, 1, -nbits);
    elsif (x=765) then return to_sfixed(0.00130718954248366004, 1, -nbits);
    elsif (x=766) then return to_sfixed(0.00130548302872062665, 1, -nbits);
    elsif (x=767) then return to_sfixed(0.00130378096479791391, 1, -nbits);
    elsif (x=768) then return to_sfixed(0.00130208333333333326, 1, -nbits);
    elsif (x=769) then return to_sfixed(0.00130039011703511056, 1, -nbits);
    elsif (x=770) then return to_sfixed(0.00129870129870129870, 1, -nbits);
    elsif (x=771) then return to_sfixed(0.00129701686121919580, 1, -nbits);
    elsif (x=772) then return to_sfixed(0.00129533678756476689, 1, -nbits);
    elsif (x=773) then return to_sfixed(0.00129366106080206996, 1, -nbits);
    elsif (x=774) then return to_sfixed(0.00129198966408268739, 1, -nbits);
    elsif (x=775) then return to_sfixed(0.00129032258064516129, 1, -nbits);
    elsif (x=776) then return to_sfixed(0.00128865979381443297, 1, -nbits);
    elsif (x=777) then return to_sfixed(0.00128700128700128696, 1, -nbits);
    elsif (x=778) then return to_sfixed(0.00128534704370179939, 1, -nbits);
    elsif (x=779) then return to_sfixed(0.00128369704749679066, 1, -nbits);
    elsif (x=780) then return to_sfixed(0.00128205128205128205, 1, -nbits);
    elsif (x=781) then return to_sfixed(0.00128040973111395642, 1, -nbits);
    elsif (x=782) then return to_sfixed(0.00127877237851662415, 1, -nbits);
    elsif (x=783) then return to_sfixed(0.00127713920817369101, 1, -nbits);
    elsif (x=784) then return to_sfixed(0.00127551020408163255, 1, -nbits);
    elsif (x=785) then return to_sfixed(0.00127388535031847127, 1, -nbits);
    elsif (x=786) then return to_sfixed(0.00127226463104325709, 1, -nbits);
    elsif (x=787) then return to_sfixed(0.00127064803049555279, 1, -nbits);
    elsif (x=788) then return to_sfixed(0.00126903553299492376, 1, -nbits);
    elsif (x=789) then return to_sfixed(0.00126742712294043085, 1, -nbits);
    elsif (x=790) then return to_sfixed(0.00126582278481012661, 1, -nbits);
    elsif (x=791) then return to_sfixed(0.00126422250316055636, 1, -nbits);
    elsif (x=792) then return to_sfixed(0.00126262626262626273, 1, -nbits);
    elsif (x=793) then return to_sfixed(0.00126103404791929382, 1, -nbits);
    elsif (x=794) then return to_sfixed(0.00125944584382871533, 1, -nbits);
    elsif (x=795) then return to_sfixed(0.00125786163522012572, 1, -nbits);
    elsif (x=796) then return to_sfixed(0.00125628140703517590, 1, -nbits);
    elsif (x=797) then return to_sfixed(0.00125470514429109150, 1, -nbits);
    elsif (x=798) then return to_sfixed(0.00125313283208020043, 1, -nbits);
    elsif (x=799) then return to_sfixed(0.00125156445556946186, 1, -nbits);
    elsif (x=800) then return to_sfixed(0.00125000000000000003, 1, -nbits);
    elsif (x=801) then return to_sfixed(0.00124843945068664171, 1, -nbits);
    elsif (x=802) then return to_sfixed(0.00124688279301745633, 1, -nbits);
    elsif (x=803) then return to_sfixed(0.00124533001245330011, 1, -nbits);
    elsif (x=804) then return to_sfixed(0.00124378109452736316, 1, -nbits);
    elsif (x=805) then return to_sfixed(0.00124223602484472054, 1, -nbits);
    elsif (x=806) then return to_sfixed(0.00124069478908188586, 1, -nbits);
    elsif (x=807) then return to_sfixed(0.00123915737298636928, 1, -nbits);
    elsif (x=808) then return to_sfixed(0.00123762376237623764, 1, -nbits);
    elsif (x=809) then return to_sfixed(0.00123609394313967851, 1, -nbits);
    elsif (x=810) then return to_sfixed(0.00123456790123456788, 1, -nbits);
    elsif (x=811) then return to_sfixed(0.00123304562268803947, 1, -nbits);
    elsif (x=812) then return to_sfixed(0.00123152709359605913, 1, -nbits);
    elsif (x=813) then return to_sfixed(0.00123001230012300127, 1, -nbits);
    elsif (x=814) then return to_sfixed(0.00122850122850122847, 1, -nbits);
    elsif (x=815) then return to_sfixed(0.00122699386503067492, 1, -nbits);
    elsif (x=816) then return to_sfixed(0.00122549019607843136, 1, -nbits);
    elsif (x=817) then return to_sfixed(0.00122399020807833527, 1, -nbits);
    elsif (x=818) then return to_sfixed(0.00122249388753056234, 1, -nbits);
    elsif (x=819) then return to_sfixed(0.00122100122100122100, 1, -nbits);
    elsif (x=820) then return to_sfixed(0.00121951219512195122, 1, -nbits);
    elsif (x=821) then return to_sfixed(0.00121802679658952490, 1, -nbits);
    elsif (x=822) then return to_sfixed(0.00121654501216545015, 1, -nbits);
    elsif (x=823) then return to_sfixed(0.00121506682867557705, 1, -nbits);
    elsif (x=824) then return to_sfixed(0.00121359223300970863, 1, -nbits);
    elsif (x=825) then return to_sfixed(0.00121212121212121212, 1, -nbits);
    elsif (x=826) then return to_sfixed(0.00121065375302663444, 1, -nbits);
    elsif (x=827) then return to_sfixed(0.00120918984280532038, 1, -nbits);
    elsif (x=828) then return to_sfixed(0.00120772946859903376, 1, -nbits);
    elsif (x=829) then return to_sfixed(0.00120627261761158014, 1, -nbits);
    elsif (x=830) then return to_sfixed(0.00120481927710843384, 1, -nbits);
    elsif (x=831) then return to_sfixed(0.00120336943441636587, 1, -nbits);
    elsif (x=832) then return to_sfixed(0.00120192307692307699, 1, -nbits);
    elsif (x=833) then return to_sfixed(0.00120048019207683065, 1, -nbits);
    elsif (x=834) then return to_sfixed(0.00119904076738609104, 1, -nbits);
    elsif (x=835) then return to_sfixed(0.00119760479041916166, 1, -nbits);
    elsif (x=836) then return to_sfixed(0.00119617224880382770, 1, -nbits);
    elsif (x=837) then return to_sfixed(0.00119474313022700112, 1, -nbits);
    elsif (x=838) then return to_sfixed(0.00119331742243436760, 1, -nbits);
    elsif (x=839) then return to_sfixed(0.00119189511323003570, 1, -nbits);
    elsif (x=840) then return to_sfixed(0.00119047619047619058, 1, -nbits);
    elsif (x=841) then return to_sfixed(0.00118906064209274662, 1, -nbits);
    elsif (x=842) then return to_sfixed(0.00118764845605700718, 1, -nbits);
    elsif (x=843) then return to_sfixed(0.00118623962040332155, 1, -nbits);
    elsif (x=844) then return to_sfixed(0.00118483412322274891, 1, -nbits);
    elsif (x=845) then return to_sfixed(0.00118343195266272191, 1, -nbits);
    elsif (x=846) then return to_sfixed(0.00118203309692671392, 1, -nbits);
    elsif (x=847) then return to_sfixed(0.00118063754427390785, 1, -nbits);
    elsif (x=848) then return to_sfixed(0.00117924528301886788, 1, -nbits);
    elsif (x=849) then return to_sfixed(0.00117785630153121310, 1, -nbits);
    elsif (x=850) then return to_sfixed(0.00117647058823529401, 1, -nbits);
    elsif (x=851) then return to_sfixed(0.00117508813160987070, 1, -nbits);
    elsif (x=852) then return to_sfixed(0.00117370892018779345, 1, -nbits);
    elsif (x=853) then return to_sfixed(0.00117233294255568573, 1, -nbits);
    elsif (x=854) then return to_sfixed(0.00117096018735362998, 1, -nbits);
    elsif (x=855) then return to_sfixed(0.00116959064327485382, 1, -nbits);
    elsif (x=856) then return to_sfixed(0.00116822429906542047, 1, -nbits);
    elsif (x=857) then return to_sfixed(0.00116686114352392055, 1, -nbits);
    elsif (x=858) then return to_sfixed(0.00116550116550116550, 1, -nbits);
    elsif (x=859) then return to_sfixed(0.00116414435389988356, 1, -nbits);
    elsif (x=860) then return to_sfixed(0.00116279069767441859, 1, -nbits);
    elsif (x=861) then return to_sfixed(0.00116144018583042973, 1, -nbits);
    elsif (x=862) then return to_sfixed(0.00116009280742459392, 1, -nbits);
    elsif (x=863) then return to_sfixed(0.00115874855156431053, 1, -nbits);
    elsif (x=864) then return to_sfixed(0.00115740740740740734, 1, -nbits);
    elsif (x=865) then return to_sfixed(0.00115606936416184978, 1, -nbits);
    elsif (x=866) then return to_sfixed(0.00115473441108545033, 1, -nbits);
    elsif (x=867) then return to_sfixed(0.00115340253748558250, 1, -nbits);
    elsif (x=868) then return to_sfixed(0.00115207373271889401, 1, -nbits);
    elsif (x=869) then return to_sfixed(0.00115074798619102417, 1, -nbits);
    elsif (x=870) then return to_sfixed(0.00114942528735632182, 1, -nbits);
    elsif (x=871) then return to_sfixed(0.00114810562571756604, 1, -nbits);
    elsif (x=872) then return to_sfixed(0.00114678899082568814, 1, -nbits);
    elsif (x=873) then return to_sfixed(0.00114547537227949604, 1, -nbits);
    elsif (x=874) then return to_sfixed(0.00114416475972540046, 1, -nbits);
    elsif (x=875) then return to_sfixed(0.00114285714285714294, 1, -nbits);
    elsif (x=876) then return to_sfixed(0.00114155251141552505, 1, -nbits);
    elsif (x=877) then return to_sfixed(0.00114025085518814143, 1, -nbits);
    elsif (x=878) then return to_sfixed(0.00113895216400911156, 1, -nbits);
    elsif (x=879) then return to_sfixed(0.00113765642775881678, 1, -nbits);
    elsif (x=880) then return to_sfixed(0.00113636363636363631, 1, -nbits);
    elsif (x=881) then return to_sfixed(0.00113507377979568669, 1, -nbits);
    elsif (x=882) then return to_sfixed(0.00113378684807256239, 1, -nbits);
    elsif (x=883) then return to_sfixed(0.00113250283125707822, 1, -nbits);
    elsif (x=884) then return to_sfixed(0.00113122171945701368, 1, -nbits);
    elsif (x=885) then return to_sfixed(0.00112994350282485880, 1, -nbits);
    elsif (x=886) then return to_sfixed(0.00112866817155756198, 1, -nbits);
    elsif (x=887) then return to_sfixed(0.00112739571589627954, 1, -nbits);
    elsif (x=888) then return to_sfixed(0.00112612612612612612, 1, -nbits);
    elsif (x=889) then return to_sfixed(0.00112485939257592812, 1, -nbits);
    elsif (x=890) then return to_sfixed(0.00112359550561797763, 1, -nbits);
    elsif (x=891) then return to_sfixed(0.00112233445566778910, 1, -nbits);
    elsif (x=892) then return to_sfixed(0.00112107623318385649, 1, -nbits);
    elsif (x=893) then return to_sfixed(0.00111982082866741322, 1, -nbits);
    elsif (x=894) then return to_sfixed(0.00111856823266219237, 1, -nbits);
    elsif (x=895) then return to_sfixed(0.00111731843575418985, 1, -nbits);
    elsif (x=896) then return to_sfixed(0.00111607142857142851, 1, -nbits);
    elsif (x=897) then return to_sfixed(0.00111482720178372350, 1, -nbits);
    elsif (x=898) then return to_sfixed(0.00111358574610244984, 1, -nbits);
    elsif (x=899) then return to_sfixed(0.00111234705228031145, 1, -nbits);
    elsif (x=900) then return to_sfixed(0.00111111111111111111, 1, -nbits);
    elsif (x=901) then return to_sfixed(0.00110987791342952277, 1, -nbits);
    elsif (x=902) then return to_sfixed(0.00110864745011086474, 1, -nbits);
    elsif (x=903) then return to_sfixed(0.00110741971207087482, 1, -nbits);
    elsif (x=904) then return to_sfixed(0.00110619469026548671, 1, -nbits);
    elsif (x=905) then return to_sfixed(0.00110497237569060782, 1, -nbits);
    elsif (x=906) then return to_sfixed(0.00110375275938189845, 1, -nbits);
    elsif (x=907) then return to_sfixed(0.00110253583241455349, 1, -nbits);
    elsif (x=908) then return to_sfixed(0.00110132158590308380, 1, -nbits);
    elsif (x=909) then return to_sfixed(0.00110011001100110005, 1, -nbits);
    elsif (x=910) then return to_sfixed(0.00109890109890109890, 1, -nbits);
    elsif (x=911) then return to_sfixed(0.00109769484083424812, 1, -nbits);
    elsif (x=912) then return to_sfixed(0.00109649122807017538, 1, -nbits);
    elsif (x=913) then return to_sfixed(0.00109529025191675792, 1, -nbits);
    elsif (x=914) then return to_sfixed(0.00109409190371991243, 1, -nbits);
    elsif (x=915) then return to_sfixed(0.00109289617486338798, 1, -nbits);
    elsif (x=916) then return to_sfixed(0.00109170305676855890, 1, -nbits);
    elsif (x=917) then return to_sfixed(0.00109051254089422033, 1, -nbits);
    elsif (x=918) then return to_sfixed(0.00108932461873638355, 1, -nbits);
    elsif (x=919) then return to_sfixed(0.00108813928182807402, 1, -nbits);
    elsif (x=920) then return to_sfixed(0.00108695652173913045, 1, -nbits);
    elsif (x=921) then return to_sfixed(0.00108577633007600439, 1, -nbits);
    elsif (x=922) then return to_sfixed(0.00108459869848156185, 1, -nbits);
    elsif (x=923) then return to_sfixed(0.00108342361863488618, 1, -nbits);
    elsif (x=924) then return to_sfixed(0.00108225108225108225, 1, -nbits);
    elsif (x=925) then return to_sfixed(0.00108108108108108110, 1, -nbits);
    elsif (x=926) then return to_sfixed(0.00107991360691144715, 1, -nbits);
    elsif (x=927) then return to_sfixed(0.00107874865156418545, 1, -nbits);
    elsif (x=928) then return to_sfixed(0.00107758620689655171, 1, -nbits);
    elsif (x=929) then return to_sfixed(0.00107642626480086104, 1, -nbits);
    elsif (x=930) then return to_sfixed(0.00107526881720430107, 1, -nbits);
    elsif (x=931) then return to_sfixed(0.00107411385606874326, 1, -nbits);
    elsif (x=932) then return to_sfixed(0.00107296137339055794, 1, -nbits);
    elsif (x=933) then return to_sfixed(0.00107181136120042871, 1, -nbits);
    elsif (x=934) then return to_sfixed(0.00107066381156316922, 1, -nbits);
    elsif (x=935) then return to_sfixed(0.00106951871657754013, 1, -nbits);
    elsif (x=936) then return to_sfixed(0.00106837606837606848, 1, -nbits);
    elsif (x=937) then return to_sfixed(0.00106723585912486666, 1, -nbits);
    elsif (x=938) then return to_sfixed(0.00106609808102345414, 1, -nbits);
    elsif (x=939) then return to_sfixed(0.00106496272630457944, 1, -nbits);
    elsif (x=940) then return to_sfixed(0.00106382978723404257, 1, -nbits);
    elsif (x=941) then return to_sfixed(0.00106269925611052066, 1, -nbits);
    elsif (x=942) then return to_sfixed(0.00106157112526539276, 1, -nbits);
    elsif (x=943) then return to_sfixed(0.00106044538706256638, 1, -nbits);
    elsif (x=944) then return to_sfixed(0.00105932203389830508, 1, -nbits);
    elsif (x=945) then return to_sfixed(0.00105820105820105827, 1, -nbits);
    elsif (x=946) then return to_sfixed(0.00105708245243128969, 1, -nbits);
    elsif (x=947) then return to_sfixed(0.00105596620908130932, 1, -nbits);
    elsif (x=948) then return to_sfixed(0.00105485232067510540, 1, -nbits);
    elsif (x=949) then return to_sfixed(0.00105374077976817695, 1, -nbits);
    elsif (x=950) then return to_sfixed(0.00105263157894736840, 1, -nbits);
    elsif (x=951) then return to_sfixed(0.00105152471083070449, 1, -nbits);
    elsif (x=952) then return to_sfixed(0.00105042016806722685, 1, -nbits);
    elsif (x=953) then return to_sfixed(0.00104931794333683109, 1, -nbits);
    elsif (x=954) then return to_sfixed(0.00104821802935010488, 1, -nbits);
    elsif (x=955) then return to_sfixed(0.00104712041884816765, 1, -nbits);
    elsif (x=956) then return to_sfixed(0.00104602510460251037, 1, -nbits);
    elsif (x=957) then return to_sfixed(0.00104493207941483814, 1, -nbits);
    elsif (x=958) then return to_sfixed(0.00104384133611691013, 1, -nbits);
    elsif (x=959) then return to_sfixed(0.00104275286757038585, 1, -nbits);
    elsif (x=960) then return to_sfixed(0.00104166666666666665, 1, -nbits);
    elsif (x=961) then return to_sfixed(0.00104058272632674307, 1, -nbits);
    elsif (x=962) then return to_sfixed(0.00103950103950103956, 1, -nbits);
    elsif (x=963) then return to_sfixed(0.00103842159916926269, 1, -nbits);
    elsif (x=964) then return to_sfixed(0.00103734439834024896, 1, -nbits);
    elsif (x=965) then return to_sfixed(0.00103626943005181342, 1, -nbits);
    elsif (x=966) then return to_sfixed(0.00103519668737060049, 1, -nbits);
    elsif (x=967) then return to_sfixed(0.00103412616339193389, 1, -nbits);
    elsif (x=968) then return to_sfixed(0.00103305785123966945, 1, -nbits);
    elsif (x=969) then return to_sfixed(0.00103199174406604739, 1, -nbits);
    elsif (x=970) then return to_sfixed(0.00103092783505154642, 1, -nbits);
    elsif (x=971) then return to_sfixed(0.00102986611740473735, 1, -nbits);
    elsif (x=972) then return to_sfixed(0.00102880658436214001, 1, -nbits);
    elsif (x=973) then return to_sfixed(0.00102774922918807813, 1, -nbits);
    elsif (x=974) then return to_sfixed(0.00102669404517453803, 1, -nbits);
    elsif (x=975) then return to_sfixed(0.00102564102564102564, 1, -nbits);
    elsif (x=976) then return to_sfixed(0.00102459016393442628, 1, -nbits);
    elsif (x=977) then return to_sfixed(0.00102354145342886389, 1, -nbits);
    elsif (x=978) then return to_sfixed(0.00102249488752556247, 1, -nbits);
    elsif (x=979) then return to_sfixed(0.00102145045965270687, 1, -nbits);
    elsif (x=980) then return to_sfixed(0.00102040816326530621, 1, -nbits);
    elsif (x=981) then return to_sfixed(0.00101936799184505615, 1, -nbits);
    elsif (x=982) then return to_sfixed(0.00101832993890020357, 1, -nbits);
    elsif (x=983) then return to_sfixed(0.00101729399796541197, 1, -nbits);
    elsif (x=984) then return to_sfixed(0.00101626016260162612, 1, -nbits);
    elsif (x=985) then return to_sfixed(0.00101522842639593914, 1, -nbits);
    elsif (x=986) then return to_sfixed(0.00101419878296146043, 1, -nbits);
    elsif (x=987) then return to_sfixed(0.00101317122593718345, 1, -nbits);
    elsif (x=988) then return to_sfixed(0.00101214574898785426, 1, -nbits);
    elsif (x=989) then return to_sfixed(0.00101112234580384231, 1, -nbits);
    elsif (x=990) then return to_sfixed(0.00101010101010101010, 1, -nbits);
    elsif (x=991) then return to_sfixed(0.00100908173562058528, 1, -nbits);
    elsif (x=992) then return to_sfixed(0.00100806451612903223, 1, -nbits);
    elsif (x=993) then return to_sfixed(0.00100704934541792548, 1, -nbits);
    elsif (x=994) then return to_sfixed(0.00100603621730382302, 1, -nbits);
    elsif (x=995) then return to_sfixed(0.00100502512562814081, 1, -nbits);
    elsif (x=996) then return to_sfixed(0.00100401606425702802, 1, -nbits);
    elsif (x=997) then return to_sfixed(0.00100300902708124373, 1, -nbits);
    elsif (x=998) then return to_sfixed(0.00100200400801603198, 1, -nbits);
    elsif (x=999) then return to_sfixed(0.00100100100100100099, 1, -nbits);
    elsif (x=1000) then return to_sfixed(0.00100000000000000002, 1, -nbits);
    elsif (x=1001) then return to_sfixed(0.00099900099900099900, 1, -nbits);
    elsif (x=1002) then return to_sfixed(0.00099800399201596798, 1, -nbits);
    elsif (x=1003) then return to_sfixed(0.00099700897308075765, 1, -nbits);
    elsif (x=1004) then return to_sfixed(0.00099601593625498006, 1, -nbits);
    elsif (x=1005) then return to_sfixed(0.00099502487562189048, 1, -nbits);
    elsif (x=1006) then return to_sfixed(0.00099403578528827028, 1, -nbits);
    elsif (x=1007) then return to_sfixed(0.00099304865938430980, 1, -nbits);
    elsif (x=1008) then return to_sfixed(0.00099206349206349201, 1, -nbits);
    elsif (x=1009) then return to_sfixed(0.00099108027750247768, 1, -nbits);
    elsif (x=1010) then return to_sfixed(0.00099009900990099011, 1, -nbits);
    elsif (x=1011) then return to_sfixed(0.00098911968348170125, 1, -nbits);
    elsif (x=1012) then return to_sfixed(0.00098814229249011851, 1, -nbits);
    elsif (x=1013) then return to_sfixed(0.00098716683119447180, 1, -nbits);
    elsif (x=1014) then return to_sfixed(0.00098619329388560163, 1, -nbits);
    elsif (x=1015) then return to_sfixed(0.00098522167487684722, 1, -nbits);
    elsif (x=1016) then return to_sfixed(0.00098425196850393699, 1, -nbits);
    elsif (x=1017) then return to_sfixed(0.00098328416912487715, 1, -nbits);
    elsif (x=1018) then return to_sfixed(0.00098231827111984276, 1, -nbits);
    elsif (x=1019) then return to_sfixed(0.00098135426889106960, 1, -nbits);
    elsif (x=1020) then return to_sfixed(0.00098039215686274508, 1, -nbits);
    elsif (x=1021) then return to_sfixed(0.00097943192948090111, 1, -nbits);
    elsif (x=1022) then return to_sfixed(0.00097847358121330719, 1, -nbits);
    elsif (x=1023) then return to_sfixed(0.00097751710654936461, 1, -nbits);
    elsif (x=1024) then return to_sfixed(0.00097656250000000000, 1, -nbits);
    elsif (x=1025) then return to_sfixed(0.00097560975609756097, 1, -nbits);
    elsif (x=1026) then return to_sfixed(0.00097465886939571145, 1, -nbits);
    elsif (x=1027) then return to_sfixed(0.00097370983446932818, 1, -nbits);
    elsif (x=1028) then return to_sfixed(0.00097276264591439690, 1, -nbits);
    elsif (x=1029) then return to_sfixed(0.00097181729834791054, 1, -nbits);
    elsif (x=1030) then return to_sfixed(0.00097087378640776695, 1, -nbits);
    elsif (x=1031) then return to_sfixed(0.00096993210475266732, 1, -nbits);
    elsif (x=1032) then return to_sfixed(0.00096899224806201549, 1, -nbits);
    elsif (x=1033) then return to_sfixed(0.00096805421103581804, 1, -nbits);
    elsif (x=1034) then return to_sfixed(0.00096711798839458415, 1, -nbits);
    elsif (x=1035) then return to_sfixed(0.00096618357487922703, 1, -nbits);
    elsif (x=1036) then return to_sfixed(0.00096525096525096527, 1, -nbits);
    elsif (x=1037) then return to_sfixed(0.00096432015429122472, 1, -nbits);
    elsif (x=1038) then return to_sfixed(0.00096339113680154141, 1, -nbits);
    elsif (x=1039) then return to_sfixed(0.00096246390760346492, 1, -nbits);
    elsif (x=1040) then return to_sfixed(0.00096153846153846159, 1, -nbits);
    elsif (x=1041) then return to_sfixed(0.00096061479346781938, 1, -nbits);
    elsif (x=1042) then return to_sfixed(0.00095969289827255275, 1, -nbits);
    elsif (x=1043) then return to_sfixed(0.00095877277085330771, 1, -nbits);
    elsif (x=1044) then return to_sfixed(0.00095785440613026815, 1, -nbits);
    elsif (x=1045) then return to_sfixed(0.00095693779904306223, 1, -nbits);
    elsif (x=1046) then return to_sfixed(0.00095602294455066918, 1, -nbits);
    elsif (x=1047) then return to_sfixed(0.00095510983763132757, 1, -nbits);
    elsif (x=1048) then return to_sfixed(0.00095419847328244271, 1, -nbits);
    elsif (x=1049) then return to_sfixed(0.00095328884652049568, 1, -nbits);
    elsif (x=1050) then return to_sfixed(0.00095238095238095238, 1, -nbits);
    elsif (x=1051) then return to_sfixed(0.00095147478591817321, 1, -nbits);
    elsif (x=1052) then return to_sfixed(0.00095057034220532319, 1, -nbits);
    elsif (x=1053) then return to_sfixed(0.00094966761633428305, 1, -nbits);
    elsif (x=1054) then return to_sfixed(0.00094876660341555979, 1, -nbits);
    elsif (x=1055) then return to_sfixed(0.00094786729857819908, 1, -nbits);
    elsif (x=1056) then return to_sfixed(0.00094696969696969700, 1, -nbits);
    elsif (x=1057) then return to_sfixed(0.00094607379375591296, 1, -nbits);
    elsif (x=1058) then return to_sfixed(0.00094517958412098301, 1, -nbits);
    elsif (x=1059) then return to_sfixed(0.00094428706326723328, 1, -nbits);
    elsif (x=1060) then return to_sfixed(0.00094339622641509435, 1, -nbits);
    elsif (x=1061) then return to_sfixed(0.00094250706880301600, 1, -nbits);
    elsif (x=1062) then return to_sfixed(0.00094161958568738226, 1, -nbits);
    elsif (x=1063) then return to_sfixed(0.00094073377234242712, 1, -nbits);
    elsif (x=1064) then return to_sfixed(0.00093984962406015032, 1, -nbits);
    elsif (x=1065) then return to_sfixed(0.00093896713615023472, 1, -nbits);
    elsif (x=1066) then return to_sfixed(0.00093808630393996248, 1, -nbits);
    elsif (x=1067) then return to_sfixed(0.00093720712277413310, 1, -nbits);
    elsif (x=1068) then return to_sfixed(0.00093632958801498128, 1, -nbits);
    elsif (x=1069) then return to_sfixed(0.00093545369504209543, 1, -nbits);
    elsif (x=1070) then return to_sfixed(0.00093457943925233649, 1, -nbits);
    elsif (x=1071) then return to_sfixed(0.00093370681605975728, 1, -nbits);
    elsif (x=1072) then return to_sfixed(0.00093283582089552237, 1, -nbits);
    elsif (x=1073) then return to_sfixed(0.00093196644920782849, 1, -nbits);
    elsif (x=1074) then return to_sfixed(0.00093109869646182495, 1, -nbits);
    elsif (x=1075) then return to_sfixed(0.00093023255813953494, 1, -nbits);
    elsif (x=1076) then return to_sfixed(0.00092936802973977691, 1, -nbits);
    elsif (x=1077) then return to_sfixed(0.00092850510677808728, 1, -nbits);
    elsif (x=1078) then return to_sfixed(0.00092764378478664194, 1, -nbits);
    elsif (x=1079) then return to_sfixed(0.00092678405931417981, 1, -nbits);
    elsif (x=1080) then return to_sfixed(0.00092592592592592596, 1, -nbits);
    elsif (x=1081) then return to_sfixed(0.00092506938020351531, 1, -nbits);
    elsif (x=1082) then return to_sfixed(0.00092421441774491681, 1, -nbits);
    elsif (x=1083) then return to_sfixed(0.00092336103416435823, 1, -nbits);
    elsif (x=1084) then return to_sfixed(0.00092250922509225090, 1, -nbits);
    elsif (x=1085) then return to_sfixed(0.00092165898617511521, 1, -nbits);
    elsif (x=1086) then return to_sfixed(0.00092081031307550648, 1, -nbits);
    elsif (x=1087) then return to_sfixed(0.00091996320147194111, 1, -nbits);
    elsif (x=1088) then return to_sfixed(0.00091911764705882352, 1, -nbits);
    elsif (x=1089) then return to_sfixed(0.00091827364554637281, 1, -nbits);
    elsif (x=1090) then return to_sfixed(0.00091743119266055051, 1, -nbits);
    elsif (x=1091) then return to_sfixed(0.00091659028414298811, 1, -nbits);
    elsif (x=1092) then return to_sfixed(0.00091575091575091575, 1, -nbits);
    elsif (x=1093) then return to_sfixed(0.00091491308325709062, 1, -nbits);
    elsif (x=1094) then return to_sfixed(0.00091407678244972577, 1, -nbits);
    elsif (x=1095) then return to_sfixed(0.00091324200913242006, 1, -nbits);
    elsif (x=1096) then return to_sfixed(0.00091240875912408756, 1, -nbits);
    elsif (x=1097) then return to_sfixed(0.00091157702825888785, 1, -nbits);
    elsif (x=1098) then return to_sfixed(0.00091074681238615665, 1, -nbits);
    elsif (x=1099) then return to_sfixed(0.00090991810737033670, 1, -nbits);
    elsif (x=1100) then return to_sfixed(0.00090909090909090909, 1, -nbits);
    elsif (x=1101) then return to_sfixed(0.00090826521344232513, 1, -nbits);
    elsif (x=1102) then return to_sfixed(0.00090744101633393826, 1, -nbits);
    elsif (x=1103) then return to_sfixed(0.00090661831368993653, 1, -nbits);
    elsif (x=1104) then return to_sfixed(0.00090579710144927537, 1, -nbits);
    elsif (x=1105) then return to_sfixed(0.00090497737556561090, 1, -nbits);
    elsif (x=1106) then return to_sfixed(0.00090415913200723324, 1, -nbits);
    elsif (x=1107) then return to_sfixed(0.00090334236675700087, 1, -nbits);
    elsif (x=1108) then return to_sfixed(0.00090252707581227440, 1, -nbits);
    elsif (x=1109) then return to_sfixed(0.00090171325518485117, 1, -nbits);
    elsif (x=1110) then return to_sfixed(0.00090090090090090091, 1, -nbits);
    elsif (x=1111) then return to_sfixed(0.00090009000900090005, 1, -nbits);
    elsif (x=1112) then return to_sfixed(0.00089928057553956839, 1, -nbits);
    elsif (x=1113) then return to_sfixed(0.00089847259658580418, 1, -nbits);
    elsif (x=1114) then return to_sfixed(0.00089766606822262122, 1, -nbits);
    elsif (x=1115) then return to_sfixed(0.00089686098654708521, 1, -nbits);
    elsif (x=1116) then return to_sfixed(0.00089605734767025090, 1, -nbits);
    elsif (x=1117) then return to_sfixed(0.00089525514771709937, 1, -nbits);
    elsif (x=1118) then return to_sfixed(0.00089445438282647585, 1, -nbits);
    elsif (x=1119) then return to_sfixed(0.00089365504915102768, 1, -nbits);
    elsif (x=1120) then return to_sfixed(0.00089285714285714283, 1, -nbits);
    elsif (x=1121) then return to_sfixed(0.00089206066012488853, 1, -nbits);
    elsif (x=1122) then return to_sfixed(0.00089126559714795004, 1, -nbits);
    elsif (x=1123) then return to_sfixed(0.00089047195013357077, 1, -nbits);
    elsif (x=1124) then return to_sfixed(0.00088967971530249106, 1, -nbits);
    elsif (x=1125) then return to_sfixed(0.00088888888888888893, 1, -nbits);
    elsif (x=1126) then return to_sfixed(0.00088809946714031975, 1, -nbits);
    elsif (x=1127) then return to_sfixed(0.00088731144631765753, 1, -nbits);
    elsif (x=1128) then return to_sfixed(0.00088652482269503544, 1, -nbits);
    elsif (x=1129) then return to_sfixed(0.00088573959255978745, 1, -nbits);
    elsif (x=1130) then return to_sfixed(0.00088495575221238937, 1, -nbits);
    elsif (x=1131) then return to_sfixed(0.00088417329796640137, 1, -nbits);
    elsif (x=1132) then return to_sfixed(0.00088339222614840988, 1, -nbits);
    elsif (x=1133) then return to_sfixed(0.00088261253309797002, 1, -nbits);
    elsif (x=1134) then return to_sfixed(0.00088183421516754845, 1, -nbits);
    elsif (x=1135) then return to_sfixed(0.00088105726872246700, 1, -nbits);
    elsif (x=1136) then return to_sfixed(0.00088028169014084509, 1, -nbits);
    elsif (x=1137) then return to_sfixed(0.00087950747581354446, 1, -nbits);
    elsif (x=1138) then return to_sfixed(0.00087873462214411243, 1, -nbits);
    elsif (x=1139) then return to_sfixed(0.00087796312554872696, 1, -nbits);
    elsif (x=1140) then return to_sfixed(0.00087719298245614037, 1, -nbits);
    elsif (x=1141) then return to_sfixed(0.00087642418930762491, 1, -nbits);
    elsif (x=1142) then return to_sfixed(0.00087565674255691769, 1, -nbits);
    elsif (x=1143) then return to_sfixed(0.00087489063867016625, 1, -nbits);
    elsif (x=1144) then return to_sfixed(0.00087412587412587413, 1, -nbits);
    elsif (x=1145) then return to_sfixed(0.00087336244541484718, 1, -nbits);
    elsif (x=1146) then return to_sfixed(0.00087260034904013963, 1, -nbits);
    elsif (x=1147) then return to_sfixed(0.00087183958151700091, 1, -nbits);
    elsif (x=1148) then return to_sfixed(0.00087108013937282230, 1, -nbits);
    elsif (x=1149) then return to_sfixed(0.00087032201914708440, 1, -nbits);
    elsif (x=1150) then return to_sfixed(0.00086956521739130438, 1, -nbits);
    elsif (x=1151) then return to_sfixed(0.00086880973066898344, 1, -nbits);
    elsif (x=1152) then return to_sfixed(0.00086805555555555551, 1, -nbits);
    elsif (x=1153) then return to_sfixed(0.00086730268863833475, 1, -nbits);
    elsif (x=1154) then return to_sfixed(0.00086655112651646442, 1, -nbits);
    elsif (x=1155) then return to_sfixed(0.00086580086580086580, 1, -nbits);
    elsif (x=1156) then return to_sfixed(0.00086505190311418688, 1, -nbits);
    elsif (x=1157) then return to_sfixed(0.00086430423509075197, 1, -nbits);
    elsif (x=1158) then return to_sfixed(0.00086355785837651119, 1, -nbits);
    elsif (x=1159) then return to_sfixed(0.00086281276962899055, 1, -nbits);
    elsif (x=1160) then return to_sfixed(0.00086206896551724137, 1, -nbits);
    elsif (x=1161) then return to_sfixed(0.00086132644272179156, 1, -nbits);
    elsif (x=1162) then return to_sfixed(0.00086058519793459555, 1, -nbits);
    elsif (x=1163) then return to_sfixed(0.00085984522785898540, 1, -nbits);
    elsif (x=1164) then return to_sfixed(0.00085910652920962198, 1, -nbits);
    elsif (x=1165) then return to_sfixed(0.00085836909871244631, 1, -nbits);
    elsif (x=1166) then return to_sfixed(0.00085763293310463120, 1, -nbits);
    elsif (x=1167) then return to_sfixed(0.00085689802913453304, 1, -nbits);
    elsif (x=1168) then return to_sfixed(0.00085616438356164379, 1, -nbits);
    elsif (x=1169) then return to_sfixed(0.00085543199315654401, 1, -nbits);
    elsif (x=1170) then return to_sfixed(0.00085470085470085470, 1, -nbits);
    elsif (x=1171) then return to_sfixed(0.00085397096498719043, 1, -nbits);
    elsif (x=1172) then return to_sfixed(0.00085324232081911264, 1, -nbits);
    elsif (x=1173) then return to_sfixed(0.00085251491901108269, 1, -nbits);
    elsif (x=1174) then return to_sfixed(0.00085178875638841568, 1, -nbits);
    elsif (x=1175) then return to_sfixed(0.00085106382978723403, 1, -nbits);
    elsif (x=1176) then return to_sfixed(0.00085034013605442174, 1, -nbits);
    elsif (x=1177) then return to_sfixed(0.00084961767204757861, 1, -nbits);
    elsif (x=1178) then return to_sfixed(0.00084889643463497452, 1, -nbits);
    elsif (x=1179) then return to_sfixed(0.00084817642069550466, 1, -nbits);
    elsif (x=1180) then return to_sfixed(0.00084745762711864404, 1, -nbits);
    elsif (x=1181) then return to_sfixed(0.00084674005080440302, 1, -nbits);
    elsif (x=1182) then return to_sfixed(0.00084602368866328254, 1, -nbits);
    elsif (x=1183) then return to_sfixed(0.00084530853761622987, 1, -nbits);
    elsif (x=1184) then return to_sfixed(0.00084459459459459464, 1, -nbits);
    elsif (x=1185) then return to_sfixed(0.00084388185654008440, 1, -nbits);
    elsif (x=1186) then return to_sfixed(0.00084317032040472171, 1, -nbits);
    elsif (x=1187) then return to_sfixed(0.00084245998315080029, 1, -nbits);
    elsif (x=1188) then return to_sfixed(0.00084175084175084171, 1, -nbits);
    elsif (x=1189) then return to_sfixed(0.00084104289318755253, 1, -nbits);
    elsif (x=1190) then return to_sfixed(0.00084033613445378156, 1, -nbits);
    elsif (x=1191) then return to_sfixed(0.00083963056255247689, 1, -nbits);
    elsif (x=1192) then return to_sfixed(0.00083892617449664428, 1, -nbits);
    elsif (x=1193) then return to_sfixed(0.00083822296730930428, 1, -nbits);
    elsif (x=1194) then return to_sfixed(0.00083752093802345060, 1, -nbits);
    elsif (x=1195) then return to_sfixed(0.00083682008368200832, 1, -nbits);
    elsif (x=1196) then return to_sfixed(0.00083612040133779263, 1, -nbits);
    elsif (x=1197) then return to_sfixed(0.00083542188805346695, 1, -nbits);
    elsif (x=1198) then return to_sfixed(0.00083472454090150253, 1, -nbits);
    elsif (x=1199) then return to_sfixed(0.00083402835696413675, 1, -nbits);
    elsif (x=1200) then return to_sfixed(0.00083333333333333339, 1, -nbits);
    elsif (x=1201) then return to_sfixed(0.00083263946711074107, 1, -nbits);
    elsif (x=1202) then return to_sfixed(0.00083194675540765393, 1, -nbits);
    elsif (x=1203) then return to_sfixed(0.00083125519534497092, 1, -nbits);
    elsif (x=1204) then return to_sfixed(0.00083056478405315617, 1, -nbits);
    elsif (x=1205) then return to_sfixed(0.00082987551867219915, 1, -nbits);
    elsif (x=1206) then return to_sfixed(0.00082918739635157548, 1, -nbits);
    elsif (x=1207) then return to_sfixed(0.00082850041425020708, 1, -nbits);
    elsif (x=1208) then return to_sfixed(0.00082781456953642384, 1, -nbits);
    elsif (x=1209) then return to_sfixed(0.00082712985938792390, 1, -nbits);
    elsif (x=1210) then return to_sfixed(0.00082644628099173552, 1, -nbits);
    elsif (x=1211) then return to_sfixed(0.00082576383154417832, 1, -nbits);
    elsif (x=1212) then return to_sfixed(0.00082508250825082509, 1, -nbits);
    elsif (x=1213) then return to_sfixed(0.00082440230832646333, 1, -nbits);
    elsif (x=1214) then return to_sfixed(0.00082372322899505767, 1, -nbits);
    elsif (x=1215) then return to_sfixed(0.00082304526748971192, 1, -nbits);
    elsif (x=1216) then return to_sfixed(0.00082236842105263153, 1, -nbits);
    elsif (x=1217) then return to_sfixed(0.00082169268693508624, 1, -nbits);
    elsif (x=1218) then return to_sfixed(0.00082101806239737272, 1, -nbits);
    elsif (x=1219) then return to_sfixed(0.00082034454470877774, 1, -nbits);
    elsif (x=1220) then return to_sfixed(0.00081967213114754098, 1, -nbits);
    elsif (x=1221) then return to_sfixed(0.00081900081900081905, 1, -nbits);
    elsif (x=1222) then return to_sfixed(0.00081833060556464816, 1, -nbits);
    elsif (x=1223) then return to_sfixed(0.00081766148814390845, 1, -nbits);
    elsif (x=1224) then return to_sfixed(0.00081699346405228761, 1, -nbits);
    elsif (x=1225) then return to_sfixed(0.00081632653061224493, 1, -nbits);
    elsif (x=1226) then return to_sfixed(0.00081566068515497557, 1, -nbits);
    elsif (x=1227) then return to_sfixed(0.00081499592502037486, 1, -nbits);
    elsif (x=1228) then return to_sfixed(0.00081433224755700329, 1, -nbits);
    elsif (x=1229) then return to_sfixed(0.00081366965012205042, 1, -nbits);
    elsif (x=1230) then return to_sfixed(0.00081300813008130081, 1, -nbits);
    elsif (x=1231) then return to_sfixed(0.00081234768480909826, 1, -nbits);
    elsif (x=1232) then return to_sfixed(0.00081168831168831174, 1, -nbits);
    elsif (x=1233) then return to_sfixed(0.00081103000811030010, 1, -nbits);
    elsif (x=1234) then return to_sfixed(0.00081037277147487841, 1, -nbits);
    elsif (x=1235) then return to_sfixed(0.00080971659919028337, 1, -nbits);
    elsif (x=1236) then return to_sfixed(0.00080906148867313920, 1, -nbits);
    elsif (x=1237) then return to_sfixed(0.00080840743734842356, 1, -nbits);
    elsif (x=1238) then return to_sfixed(0.00080775444264943462, 1, -nbits);
    elsif (x=1239) then return to_sfixed(0.00080710250201775622, 1, -nbits);
    elsif (x=1240) then return to_sfixed(0.00080645161290322581, 1, -nbits);
    elsif (x=1241) then return to_sfixed(0.00080580177276390005, 1, -nbits);
    elsif (x=1242) then return to_sfixed(0.00080515297906602254, 1, -nbits);
    elsif (x=1243) then return to_sfixed(0.00080450522928399030, 1, -nbits);
    elsif (x=1244) then return to_sfixed(0.00080385852090032153, 1, -nbits);
    elsif (x=1245) then return to_sfixed(0.00080321285140562252, 1, -nbits);
    elsif (x=1246) then return to_sfixed(0.00080256821829855537, 1, -nbits);
    elsif (x=1247) then return to_sfixed(0.00080192461908580592, 1, -nbits);
    elsif (x=1248) then return to_sfixed(0.00080128205128205125, 1, -nbits);
    elsif (x=1249) then return to_sfixed(0.00080064051240992789, 1, -nbits);
    elsif (x=1250) then return to_sfixed(0.00080000000000000004, 1, -nbits);
    elsif (x=1251) then return to_sfixed(0.00079936051159072740, 1, -nbits);
    elsif (x=1252) then return to_sfixed(0.00079872204472843447, 1, -nbits);
    elsif (x=1253) then return to_sfixed(0.00079808459696727857, 1, -nbits);
    elsif (x=1254) then return to_sfixed(0.00079744816586921851, 1, -nbits);
    elsif (x=1255) then return to_sfixed(0.00079681274900398409, 1, -nbits);
    elsif (x=1256) then return to_sfixed(0.00079617834394904463, 1, -nbits);
    elsif (x=1257) then return to_sfixed(0.00079554494828957840, 1, -nbits);
    elsif (x=1258) then return to_sfixed(0.00079491255961844202, 1, -nbits);
    elsif (x=1259) then return to_sfixed(0.00079428117553613975, 1, -nbits);
    elsif (x=1260) then return to_sfixed(0.00079365079365079365, 1, -nbits);
    elsif (x=1261) then return to_sfixed(0.00079302141157811261, 1, -nbits);
    elsif (x=1262) then return to_sfixed(0.00079239302694136295, 1, -nbits);
    elsif (x=1263) then return to_sfixed(0.00079176563737133805, 1, -nbits);
    elsif (x=1264) then return to_sfixed(0.00079113924050632910, 1, -nbits);
    elsif (x=1265) then return to_sfixed(0.00079051383399209485, 1, -nbits);
    elsif (x=1266) then return to_sfixed(0.00078988941548183253, 1, -nbits);
    elsif (x=1267) then return to_sfixed(0.00078926598263614838, 1, -nbits);
    elsif (x=1268) then return to_sfixed(0.00078864353312302837, 1, -nbits);
    elsif (x=1269) then return to_sfixed(0.00078802206461780935, 1, -nbits);
    elsif (x=1270) then return to_sfixed(0.00078740157480314960, 1, -nbits);
    elsif (x=1271) then return to_sfixed(0.00078678206136900079, 1, -nbits);
    elsif (x=1272) then return to_sfixed(0.00078616352201257866, 1, -nbits);
    elsif (x=1273) then return to_sfixed(0.00078554595443833470, 1, -nbits);
    elsif (x=1274) then return to_sfixed(0.00078492935635792783, 1, -nbits);
    elsif (x=1275) then return to_sfixed(0.00078431372549019605, 1, -nbits);
    elsif (x=1276) then return to_sfixed(0.00078369905956112850, 1, -nbits);
    elsif (x=1277) then return to_sfixed(0.00078308535630383712, 1, -nbits);
    elsif (x=1278) then return to_sfixed(0.00078247261345852897, 1, -nbits);
    elsif (x=1279) then return to_sfixed(0.00078186082877247849, 1, -nbits);
    elsif (x=1280) then return to_sfixed(0.00078125000000000004, 1, -nbits);
    elsif (x=1281) then return to_sfixed(0.00078064012490241998, 1, -nbits);
    elsif (x=1282) then return to_sfixed(0.00078003120124804995, 1, -nbits);
    elsif (x=1283) then return to_sfixed(0.00077942322681215901, 1, -nbits);
    elsif (x=1284) then return to_sfixed(0.00077881619937694702, 1, -nbits);
    elsif (x=1285) then return to_sfixed(0.00077821011673151756, 1, -nbits);
    elsif (x=1286) then return to_sfixed(0.00077760497667185070, 1, -nbits);
    elsif (x=1287) then return to_sfixed(0.00077700077700077700, 1, -nbits);
    elsif (x=1288) then return to_sfixed(0.00077639751552795026, 1, -nbits);
    elsif (x=1289) then return to_sfixed(0.00077579519006982156, 1, -nbits);
    elsif (x=1290) then return to_sfixed(0.00077519379844961239, 1, -nbits);
    elsif (x=1291) then return to_sfixed(0.00077459333849728897, 1, -nbits);
    elsif (x=1292) then return to_sfixed(0.00077399380804953565, 1, -nbits);
    elsif (x=1293) then return to_sfixed(0.00077339520494972935, 1, -nbits);
    elsif (x=1294) then return to_sfixed(0.00077279752704791343, 1, -nbits);
    elsif (x=1295) then return to_sfixed(0.00077220077220077220, 1, -nbits);
    elsif (x=1296) then return to_sfixed(0.00077160493827160490, 1, -nbits);
    elsif (x=1297) then return to_sfixed(0.00077101002313030066, 1, -nbits);
    elsif (x=1298) then return to_sfixed(0.00077041602465331282, 1, -nbits);
    elsif (x=1299) then return to_sfixed(0.00076982294072363352, 1, -nbits);
    elsif (x=1300) then return to_sfixed(0.00076923076923076923, 1, -nbits);
    elsif (x=1301) then return to_sfixed(0.00076863950807071484, 1, -nbits);
    elsif (x=1302) then return to_sfixed(0.00076804915514592934, 1, -nbits);
    elsif (x=1303) then return to_sfixed(0.00076745970836531081, 1, -nbits);
    elsif (x=1304) then return to_sfixed(0.00076687116564417180, 1, -nbits);
    elsif (x=1305) then return to_sfixed(0.00076628352490421458, 1, -nbits);
    elsif (x=1306) then return to_sfixed(0.00076569678407350692, 1, -nbits);
    elsif (x=1307) then return to_sfixed(0.00076511094108645751, 1, -nbits);
    elsif (x=1308) then return to_sfixed(0.00076452599388379206, 1, -nbits);
    elsif (x=1309) then return to_sfixed(0.00076394194041252863, 1, -nbits);
    elsif (x=1310) then return to_sfixed(0.00076335877862595419, 1, -nbits);
    elsif (x=1311) then return to_sfixed(0.00076277650648360034, 1, -nbits);
    elsif (x=1312) then return to_sfixed(0.00076219512195121954, 1, -nbits);
    elsif (x=1313) then return to_sfixed(0.00076161462300076163, 1, -nbits);
    elsif (x=1314) then return to_sfixed(0.00076103500761035003, 1, -nbits);
    elsif (x=1315) then return to_sfixed(0.00076045627376425851, 1, -nbits);
    elsif (x=1316) then return to_sfixed(0.00075987841945288754, 1, -nbits);
    elsif (x=1317) then return to_sfixed(0.00075930144267274111, 1, -nbits);
    elsif (x=1318) then return to_sfixed(0.00075872534142640367, 1, -nbits);
    elsif (x=1319) then return to_sfixed(0.00075815011372251705, 1, -nbits);
    elsif (x=1320) then return to_sfixed(0.00075757575757575758, 1, -nbits);
    elsif (x=1321) then return to_sfixed(0.00075700227100681302, 1, -nbits);
    elsif (x=1322) then return to_sfixed(0.00075642965204236008, 1, -nbits);
    elsif (x=1323) then return to_sfixed(0.00075585789871504159, 1, -nbits);
    elsif (x=1324) then return to_sfixed(0.00075528700906344411, 1, -nbits);
    elsif (x=1325) then return to_sfixed(0.00075471698113207543, 1, -nbits);
    elsif (x=1326) then return to_sfixed(0.00075414781297134241, 1, -nbits);
    elsif (x=1327) then return to_sfixed(0.00075357950263752827, 1, -nbits);
    elsif (x=1328) then return to_sfixed(0.00075301204819277112, 1, -nbits);
    elsif (x=1329) then return to_sfixed(0.00075244544770504136, 1, -nbits);
    elsif (x=1330) then return to_sfixed(0.00075187969924812035, 1, -nbits);
    elsif (x=1331) then return to_sfixed(0.00075131480090157780, 1, -nbits);
    elsif (x=1332) then return to_sfixed(0.00075075075075075074, 1, -nbits);
    elsif (x=1333) then return to_sfixed(0.00075018754688672170, 1, -nbits);
    elsif (x=1334) then return to_sfixed(0.00074962518740629683, 1, -nbits);
    elsif (x=1335) then return to_sfixed(0.00074906367041198505, 1, -nbits);
    elsif (x=1336) then return to_sfixed(0.00074850299401197609, 1, -nbits);
    elsif (x=1337) then return to_sfixed(0.00074794315632011965, 1, -nbits);
    elsif (x=1338) then return to_sfixed(0.00074738415545590436, 1, -nbits);
    elsif (x=1339) then return to_sfixed(0.00074682598954443620, 1, -nbits);
    elsif (x=1340) then return to_sfixed(0.00074626865671641792, 1, -nbits);
    elsif (x=1341) then return to_sfixed(0.00074571215510812821, 1, -nbits);
    elsif (x=1342) then return to_sfixed(0.00074515648286140089, 1, -nbits);
    elsif (x=1343) then return to_sfixed(0.00074460163812360388, 1, -nbits);
    elsif (x=1344) then return to_sfixed(0.00074404761904761901, 1, -nbits);
    elsif (x=1345) then return to_sfixed(0.00074349442379182155, 1, -nbits);
    elsif (x=1346) then return to_sfixed(0.00074294205052005940, 1, -nbits);
    elsif (x=1347) then return to_sfixed(0.00074239049740163323, 1, -nbits);
    elsif (x=1348) then return to_sfixed(0.00074183976261127599, 1, -nbits);
    elsif (x=1349) then return to_sfixed(0.00074128984432913266, 1, -nbits);
    elsif (x=1350) then return to_sfixed(0.00074074074074074070, 1, -nbits);
    elsif (x=1351) then return to_sfixed(0.00074019245003700959, 1, -nbits);
    elsif (x=1352) then return to_sfixed(0.00073964497041420117, 1, -nbits);
    elsif (x=1353) then return to_sfixed(0.00073909830007390983, 1, -nbits);
    elsif (x=1354) then return to_sfixed(0.00073855243722304289, 1, -nbits);
    elsif (x=1355) then return to_sfixed(0.00073800738007380072, 1, -nbits);
    elsif (x=1356) then return to_sfixed(0.00073746312684365781, 1, -nbits);
    elsif (x=1357) then return to_sfixed(0.00073691967575534268, 1, -nbits);
    elsif (x=1358) then return to_sfixed(0.00073637702503681884, 1, -nbits);
    elsif (x=1359) then return to_sfixed(0.00073583517292126564, 1, -nbits);
    elsif (x=1360) then return to_sfixed(0.00073529411764705881, 1, -nbits);
    elsif (x=1361) then return to_sfixed(0.00073475385745775160, 1, -nbits);
    elsif (x=1362) then return to_sfixed(0.00073421439060205576, 1, -nbits);
    elsif (x=1363) then return to_sfixed(0.00073367571533382249, 1, -nbits);
    elsif (x=1364) then return to_sfixed(0.00073313782991202346, 1, -nbits);
    elsif (x=1365) then return to_sfixed(0.00073260073260073260, 1, -nbits);
    elsif (x=1366) then return to_sfixed(0.00073206442166910690, 1, -nbits);
    elsif (x=1367) then return to_sfixed(0.00073152889539136799, 1, -nbits);
    elsif (x=1368) then return to_sfixed(0.00073099415204678359, 1, -nbits);
    elsif (x=1369) then return to_sfixed(0.00073046018991964939, 1, -nbits);
    elsif (x=1370) then return to_sfixed(0.00072992700729927003, 1, -nbits);
    elsif (x=1371) then return to_sfixed(0.00072939460247994166, 1, -nbits);
    elsif (x=1372) then return to_sfixed(0.00072886297376093293, 1, -nbits);
    elsif (x=1373) then return to_sfixed(0.00072833211944646763, 1, -nbits);
    elsif (x=1374) then return to_sfixed(0.00072780203784570600, 1, -nbits);
    elsif (x=1375) then return to_sfixed(0.00072727272727272723, 1, -nbits);
    elsif (x=1376) then return to_sfixed(0.00072674418604651162, 1, -nbits);
    elsif (x=1377) then return to_sfixed(0.00072621641249092229, 1, -nbits);
    elsif (x=1378) then return to_sfixed(0.00072568940493468795, 1, -nbits);
    elsif (x=1379) then return to_sfixed(0.00072516316171138508, 1, -nbits);
    elsif (x=1380) then return to_sfixed(0.00072463768115942030, 1, -nbits);
    elsif (x=1381) then return to_sfixed(0.00072411296162201298, 1, -nbits);
    elsif (x=1382) then return to_sfixed(0.00072358900144717795, 1, -nbits);
    elsif (x=1383) then return to_sfixed(0.00072306579898770787, 1, -nbits);
    elsif (x=1384) then return to_sfixed(0.00072254335260115603, 1, -nbits);
    elsif (x=1385) then return to_sfixed(0.00072202166064981946, 1, -nbits);
    elsif (x=1386) then return to_sfixed(0.00072150072150072150, 1, -nbits);
    elsif (x=1387) then return to_sfixed(0.00072098053352559477, 1, -nbits);
    elsif (x=1388) then return to_sfixed(0.00072046109510086451, 1, -nbits);
    elsif (x=1389) then return to_sfixed(0.00071994240460763136, 1, -nbits);
    elsif (x=1390) then return to_sfixed(0.00071942446043165469, 1, -nbits);
    elsif (x=1391) then return to_sfixed(0.00071890726096333576, 1, -nbits);
    elsif (x=1392) then return to_sfixed(0.00071839080459770114, 1, -nbits);
    elsif (x=1393) then return to_sfixed(0.00071787508973438624, 1, -nbits);
    elsif (x=1394) then return to_sfixed(0.00071736011477761840, 1, -nbits);
    elsif (x=1395) then return to_sfixed(0.00071684587813620072, 1, -nbits);
    elsif (x=1396) then return to_sfixed(0.00071633237822349568, 1, -nbits);
    elsif (x=1397) then return to_sfixed(0.00071581961345740870, 1, -nbits);
    elsif (x=1398) then return to_sfixed(0.00071530758226037196, 1, -nbits);
    elsif (x=1399) then return to_sfixed(0.00071479628305932811, 1, -nbits);
    elsif (x=1400) then return to_sfixed(0.00071428571428571429, 1, -nbits);
    elsif (x=1401) then return to_sfixed(0.00071377587437544611, 1, -nbits);
    elsif (x=1402) then return to_sfixed(0.00071326676176890159, 1, -nbits);
    elsif (x=1403) then return to_sfixed(0.00071275837491090524, 1, -nbits);
    elsif (x=1404) then return to_sfixed(0.00071225071225071229, 1, -nbits);
    elsif (x=1405) then return to_sfixed(0.00071174377224199293, 1, -nbits);
    elsif (x=1406) then return to_sfixed(0.00071123755334281653, 1, -nbits);
    elsif (x=1407) then return to_sfixed(0.00071073205401563609, 1, -nbits);
    elsif (x=1408) then return to_sfixed(0.00071022727272727275, 1, -nbits);
    elsif (x=1409) then return to_sfixed(0.00070972320794889996, 1, -nbits);
    elsif (x=1410) then return to_sfixed(0.00070921985815602842, 1, -nbits);
    elsif (x=1411) then return to_sfixed(0.00070871722182849046, 1, -nbits);
    elsif (x=1412) then return to_sfixed(0.00070821529745042496, 1, -nbits);
    elsif (x=1413) then return to_sfixed(0.00070771408351026188, 1, -nbits);
    elsif (x=1414) then return to_sfixed(0.00070721357850070724, 1, -nbits);
    elsif (x=1415) then return to_sfixed(0.00070671378091872788, 1, -nbits);
    elsif (x=1416) then return to_sfixed(0.00070621468926553672, 1, -nbits);
    elsif (x=1417) then return to_sfixed(0.00070571630204657732, 1, -nbits);
    elsif (x=1418) then return to_sfixed(0.00070521861777150916, 1, -nbits);
    elsif (x=1419) then return to_sfixed(0.00070472163495419312, 1, -nbits);
    elsif (x=1420) then return to_sfixed(0.00070422535211267609, 1, -nbits);
    elsif (x=1421) then return to_sfixed(0.00070372976776917663, 1, -nbits);
    elsif (x=1422) then return to_sfixed(0.00070323488045007034, 1, -nbits);
    elsif (x=1423) then return to_sfixed(0.00070274068868587491, 1, -nbits);
    elsif (x=1424) then return to_sfixed(0.00070224719101123594, 1, -nbits);
    elsif (x=1425) then return to_sfixed(0.00070175438596491223, 1, -nbits);
    elsif (x=1426) then return to_sfixed(0.00070126227208976155, 1, -nbits);
    elsif (x=1427) then return to_sfixed(0.00070077084793272596, 1, -nbits);
    elsif (x=1428) then return to_sfixed(0.00070028011204481793, 1, -nbits);
    elsif (x=1429) then return to_sfixed(0.00069979006298110562, 1, -nbits);
    elsif (x=1430) then return to_sfixed(0.00069930069930069930, 1, -nbits);
    elsif (x=1431) then return to_sfixed(0.00069881201956673651, 1, -nbits);
    elsif (x=1432) then return to_sfixed(0.00069832402234636874, 1, -nbits);
    elsif (x=1433) then return to_sfixed(0.00069783670621074664, 1, -nbits);
    elsif (x=1434) then return to_sfixed(0.00069735006973500695, 1, -nbits);
    elsif (x=1435) then return to_sfixed(0.00069686411149825784, 1, -nbits);
    elsif (x=1436) then return to_sfixed(0.00069637883008356546, 1, -nbits);
    elsif (x=1437) then return to_sfixed(0.00069589422407794019, 1, -nbits);
    elsif (x=1438) then return to_sfixed(0.00069541029207232264, 1, -nbits);
    elsif (x=1439) then return to_sfixed(0.00069492703266157052, 1, -nbits);
    elsif (x=1440) then return to_sfixed(0.00069444444444444447, 1, -nbits);
    elsif (x=1441) then return to_sfixed(0.00069396252602359470, 1, -nbits);
    elsif (x=1442) then return to_sfixed(0.00069348127600554787, 1, -nbits);
    elsif (x=1443) then return to_sfixed(0.00069300069300069300, 1, -nbits);
    elsif (x=1444) then return to_sfixed(0.00069252077562326870, 1, -nbits);
    elsif (x=1445) then return to_sfixed(0.00069204152249134946, 1, -nbits);
    elsif (x=1446) then return to_sfixed(0.00069156293222683268, 1, -nbits);
    elsif (x=1447) then return to_sfixed(0.00069108500345542499, 1, -nbits);
    elsif (x=1448) then return to_sfixed(0.00069060773480662981, 1, -nbits);
    elsif (x=1449) then return to_sfixed(0.00069013112491373362, 1, -nbits);
    elsif (x=1450) then return to_sfixed(0.00068965517241379305, 1, -nbits);
    elsif (x=1451) then return to_sfixed(0.00068917987594762232, 1, -nbits);
    elsif (x=1452) then return to_sfixed(0.00068870523415977963, 1, -nbits);
    elsif (x=1453) then return to_sfixed(0.00068823124569855469, 1, -nbits);
    elsif (x=1454) then return to_sfixed(0.00068775790921595599, 1, -nbits);
    elsif (x=1455) then return to_sfixed(0.00068728522336769765, 1, -nbits);
    elsif (x=1456) then return to_sfixed(0.00068681318681318687, 1, -nbits);
    elsif (x=1457) then return to_sfixed(0.00068634179821551130, 1, -nbits);
    elsif (x=1458) then return to_sfixed(0.00068587105624142656, 1, -nbits);
    elsif (x=1459) then return to_sfixed(0.00068540095956134343, 1, -nbits);
    elsif (x=1460) then return to_sfixed(0.00068493150684931507, 1, -nbits);
    elsif (x=1461) then return to_sfixed(0.00068446269678302531, 1, -nbits);
    elsif (x=1462) then return to_sfixed(0.00068399452804377564, 1, -nbits);
    elsif (x=1463) then return to_sfixed(0.00068352699931647305, 1, -nbits);
    elsif (x=1464) then return to_sfixed(0.00068306010928961749, 1, -nbits);
    elsif (x=1465) then return to_sfixed(0.00068259385665529011, 1, -nbits);
    elsif (x=1466) then return to_sfixed(0.00068212824010914052, 1, -nbits);
    elsif (x=1467) then return to_sfixed(0.00068166325835037494, 1, -nbits);
    elsif (x=1468) then return to_sfixed(0.00068119891008174384, 1, -nbits);
    elsif (x=1469) then return to_sfixed(0.00068073519400953025, 1, -nbits);
    elsif (x=1470) then return to_sfixed(0.00068027210884353737, 1, -nbits);
    elsif (x=1471) then return to_sfixed(0.00067980965329707678, 1, -nbits);
    elsif (x=1472) then return to_sfixed(0.00067934782608695650, 1, -nbits);
    elsif (x=1473) then return to_sfixed(0.00067888662593346908, 1, -nbits);
    elsif (x=1474) then return to_sfixed(0.00067842605156037987, 1, -nbits);
    elsif (x=1475) then return to_sfixed(0.00067796610169491530, 1, -nbits);
    elsif (x=1476) then return to_sfixed(0.00067750677506775068, 1, -nbits);
    elsif (x=1477) then return to_sfixed(0.00067704807041299930, 1, -nbits);
    elsif (x=1478) then return to_sfixed(0.00067658998646820032, 1, -nbits);
    elsif (x=1479) then return to_sfixed(0.00067613252197430695, 1, -nbits);
    elsif (x=1480) then return to_sfixed(0.00067567567567567571, 1, -nbits);
    elsif (x=1481) then return to_sfixed(0.00067521944632005406, 1, -nbits);
    elsif (x=1482) then return to_sfixed(0.00067476383265856947, 1, -nbits);
    elsif (x=1483) then return to_sfixed(0.00067430883344571813, 1, -nbits);
    elsif (x=1484) then return to_sfixed(0.00067385444743935314, 1, -nbits);
    elsif (x=1485) then return to_sfixed(0.00067340067340067344, 1, -nbits);
    elsif (x=1486) then return to_sfixed(0.00067294751009421266, 1, -nbits);
    elsif (x=1487) then return to_sfixed(0.00067249495628782783, 1, -nbits);
    elsif (x=1488) then return to_sfixed(0.00067204301075268823, 1, -nbits);
    elsif (x=1489) then return to_sfixed(0.00067159167226326397, 1, -nbits);
    elsif (x=1490) then return to_sfixed(0.00067114093959731540, 1, -nbits);
    elsif (x=1491) then return to_sfixed(0.00067069081153588194, 1, -nbits);
    elsif (x=1492) then return to_sfixed(0.00067024128686327079, 1, -nbits);
    elsif (x=1493) then return to_sfixed(0.00066979236436704619, 1, -nbits);
    elsif (x=1494) then return to_sfixed(0.00066934404283801872, 1, -nbits);
    elsif (x=1495) then return to_sfixed(0.00066889632107023408, 1, -nbits);
    elsif (x=1496) then return to_sfixed(0.00066844919786096253, 1, -nbits);
    elsif (x=1497) then return to_sfixed(0.00066800267201068810, 1, -nbits);
    elsif (x=1498) then return to_sfixed(0.00066755674232309744, 1, -nbits);
    elsif (x=1499) then return to_sfixed(0.00066711140760506999, 1, -nbits);
    elsif (x=1500) then return to_sfixed(0.00066666666666666664, 1, -nbits);
    elsif (x=1501) then return to_sfixed(0.00066622251832111927, 1, -nbits);
    elsif (x=1502) then return to_sfixed(0.00066577896138482028, 1, -nbits);
    elsif (x=1503) then return to_sfixed(0.00066533599467731206, 1, -nbits);
    elsif (x=1504) then return to_sfixed(0.00066489361702127658, 1, -nbits);
    elsif (x=1505) then return to_sfixed(0.00066445182724252495, 1, -nbits);
    elsif (x=1506) then return to_sfixed(0.00066401062416998667, 1, -nbits);
    elsif (x=1507) then return to_sfixed(0.00066357000663570006, 1, -nbits);
    elsif (x=1508) then return to_sfixed(0.00066312997347480103, 1, -nbits);
    elsif (x=1509) then return to_sfixed(0.00066269052352551359, 1, -nbits);
    elsif (x=1510) then return to_sfixed(0.00066225165562913907, 1, -nbits);
    elsif (x=1511) then return to_sfixed(0.00066181336863004633, 1, -nbits);
    elsif (x=1512) then return to_sfixed(0.00066137566137566134, 1, -nbits);
    elsif (x=1513) then return to_sfixed(0.00066093853271645734, 1, -nbits);
    elsif (x=1514) then return to_sfixed(0.00066050198150594452, 1, -nbits);
    elsif (x=1515) then return to_sfixed(0.00066006600660066007, 1, -nbits);
    elsif (x=1516) then return to_sfixed(0.00065963060686015829, 1, -nbits);
    elsif (x=1517) then return to_sfixed(0.00065919578114700061, 1, -nbits);
    elsif (x=1518) then return to_sfixed(0.00065876152832674575, 1, -nbits);
    elsif (x=1519) then return to_sfixed(0.00065832784726793940, 1, -nbits);
    elsif (x=1520) then return to_sfixed(0.00065789473684210525, 1, -nbits);
    elsif (x=1521) then return to_sfixed(0.00065746219592373442, 1, -nbits);
    elsif (x=1522) then return to_sfixed(0.00065703022339027597, 1, -nbits);
    elsif (x=1523) then return to_sfixed(0.00065659881812212733, 1, -nbits);
    elsif (x=1524) then return to_sfixed(0.00065616797900262466, 1, -nbits);
    elsif (x=1525) then return to_sfixed(0.00065573770491803279, 1, -nbits);
    elsif (x=1526) then return to_sfixed(0.00065530799475753605, 1, -nbits);
    elsif (x=1527) then return to_sfixed(0.00065487884741322858, 1, -nbits);
    elsif (x=1528) then return to_sfixed(0.00065445026178010475, 1, -nbits);
    elsif (x=1529) then return to_sfixed(0.00065402223675604975, 1, -nbits);
    elsif (x=1530) then return to_sfixed(0.00065359477124183002, 1, -nbits);
    elsif (x=1531) then return to_sfixed(0.00065316786414108428, 1, -nbits);
    elsif (x=1532) then return to_sfixed(0.00065274151436031332, 1, -nbits);
    elsif (x=1533) then return to_sfixed(0.00065231572080887146, 1, -nbits);
    elsif (x=1534) then return to_sfixed(0.00065189048239895696, 1, -nbits);
    elsif (x=1535) then return to_sfixed(0.00065146579804560263, 1, -nbits);
    elsif (x=1536) then return to_sfixed(0.00065104166666666663, 1, -nbits);
    elsif (x=1537) then return to_sfixed(0.00065061808718282373, 1, -nbits);
    elsif (x=1538) then return to_sfixed(0.00065019505851755528, 1, -nbits);
    elsif (x=1539) then return to_sfixed(0.00064977257959714096, 1, -nbits);
    elsif (x=1540) then return to_sfixed(0.00064935064935064935, 1, -nbits);
    elsif (x=1541) then return to_sfixed(0.00064892926670992858, 1, -nbits);
    elsif (x=1542) then return to_sfixed(0.00064850843060959790, 1, -nbits);
    elsif (x=1543) then return to_sfixed(0.00064808813998703824, 1, -nbits);
    elsif (x=1544) then return to_sfixed(0.00064766839378238344, 1, -nbits);
    elsif (x=1545) then return to_sfixed(0.00064724919093851134, 1, -nbits);
    elsif (x=1546) then return to_sfixed(0.00064683053040103498, 1, -nbits);
    elsif (x=1547) then return to_sfixed(0.00064641241111829345, 1, -nbits);
    elsif (x=1548) then return to_sfixed(0.00064599483204134370, 1, -nbits);
    elsif (x=1549) then return to_sfixed(0.00064557779212395089, 1, -nbits);
    elsif (x=1550) then return to_sfixed(0.00064516129032258064, 1, -nbits);
    elsif (x=1551) then return to_sfixed(0.00064474532559638943, 1, -nbits);
    elsif (x=1552) then return to_sfixed(0.00064432989690721648, 1, -nbits);
    elsif (x=1553) then return to_sfixed(0.00064391500321957500, 1, -nbits);
    elsif (x=1554) then return to_sfixed(0.00064350064350064348, 1, -nbits);
    elsif (x=1555) then return to_sfixed(0.00064308681672025725, 1, -nbits);
    elsif (x=1556) then return to_sfixed(0.00064267352185089970, 1, -nbits);
    elsif (x=1557) then return to_sfixed(0.00064226075786769424, 1, -nbits);
    elsif (x=1558) then return to_sfixed(0.00064184852374839533, 1, -nbits);
    elsif (x=1559) then return to_sfixed(0.00064143681847338033, 1, -nbits);
    elsif (x=1560) then return to_sfixed(0.00064102564102564103, 1, -nbits);
    elsif (x=1561) then return to_sfixed(0.00064061499039077510, 1, -nbits);
    elsif (x=1562) then return to_sfixed(0.00064020486555697821, 1, -nbits);
    elsif (x=1563) then return to_sfixed(0.00063979526551503517, 1, -nbits);
    elsif (x=1564) then return to_sfixed(0.00063938618925831207, 1, -nbits);
    elsif (x=1565) then return to_sfixed(0.00063897763578274762, 1, -nbits);
    elsif (x=1566) then return to_sfixed(0.00063856960408684551, 1, -nbits);
    elsif (x=1567) then return to_sfixed(0.00063816209317166565, 1, -nbits);
    elsif (x=1568) then return to_sfixed(0.00063775510204081628, 1, -nbits);
    elsif (x=1569) then return to_sfixed(0.00063734862970044612, 1, -nbits);
    elsif (x=1570) then return to_sfixed(0.00063694267515923564, 1, -nbits);
    elsif (x=1571) then return to_sfixed(0.00063653723742838951, 1, -nbits);
    elsif (x=1572) then return to_sfixed(0.00063613231552162855, 1, -nbits);
    elsif (x=1573) then return to_sfixed(0.00063572790845518119, 1, -nbits);
    elsif (x=1574) then return to_sfixed(0.00063532401524777639, 1, -nbits);
    elsif (x=1575) then return to_sfixed(0.00063492063492063492, 1, -nbits);
    elsif (x=1576) then return to_sfixed(0.00063451776649746188, 1, -nbits);
    elsif (x=1577) then return to_sfixed(0.00063411540900443881, 1, -nbits);
    elsif (x=1578) then return to_sfixed(0.00063371356147021542, 1, -nbits);
    elsif (x=1579) then return to_sfixed(0.00063331222292590248, 1, -nbits);
    elsif (x=1580) then return to_sfixed(0.00063291139240506330, 1, -nbits);
    elsif (x=1581) then return to_sfixed(0.00063251106894370653, 1, -nbits);
    elsif (x=1582) then return to_sfixed(0.00063211125158027818, 1, -nbits);
    elsif (x=1583) then return to_sfixed(0.00063171193935565378, 1, -nbits);
    elsif (x=1584) then return to_sfixed(0.00063131313131313137, 1, -nbits);
    elsif (x=1585) then return to_sfixed(0.00063091482649842276, 1, -nbits);
    elsif (x=1586) then return to_sfixed(0.00063051702395964691, 1, -nbits);
    elsif (x=1587) then return to_sfixed(0.00063011972274732201, 1, -nbits);
    elsif (x=1588) then return to_sfixed(0.00062972292191435767, 1, -nbits);
    elsif (x=1589) then return to_sfixed(0.00062932662051604787, 1, -nbits);
    elsif (x=1590) then return to_sfixed(0.00062893081761006286, 1, -nbits);
    elsif (x=1591) then return to_sfixed(0.00062853551225644250, 1, -nbits);
    elsif (x=1592) then return to_sfixed(0.00062814070351758795, 1, -nbits);
    elsif (x=1593) then return to_sfixed(0.00062774639045825491, 1, -nbits);
    elsif (x=1594) then return to_sfixed(0.00062735257214554575, 1, -nbits);
    elsif (x=1595) then return to_sfixed(0.00062695924764890286, 1, -nbits);
    elsif (x=1596) then return to_sfixed(0.00062656641604010022, 1, -nbits);
    elsif (x=1597) then return to_sfixed(0.00062617407639323729, 1, -nbits);
    elsif (x=1598) then return to_sfixed(0.00062578222778473093, 1, -nbits);
    elsif (x=1599) then return to_sfixed(0.00062539086929330832, 1, -nbits);
    elsif (x=1600) then return to_sfixed(0.00062500000000000001, 1, -nbits);
    elsif (x=1601) then return to_sfixed(0.00062460961898813238, 1, -nbits);
    elsif (x=1602) then return to_sfixed(0.00062421972534332086, 1, -nbits);
    elsif (x=1603) then return to_sfixed(0.00062383031815346226, 1, -nbits);
    elsif (x=1604) then return to_sfixed(0.00062344139650872816, 1, -nbits);
    elsif (x=1605) then return to_sfixed(0.00062305295950155766, 1, -nbits);
    elsif (x=1606) then return to_sfixed(0.00062266500622665006, 1, -nbits);
    elsif (x=1607) then return to_sfixed(0.00062227753578095830, 1, -nbits);
    elsif (x=1608) then return to_sfixed(0.00062189054726368158, 1, -nbits);
    elsif (x=1609) then return to_sfixed(0.00062150403977625850, 1, -nbits);
    elsif (x=1610) then return to_sfixed(0.00062111801242236027, 1, -nbits);
    elsif (x=1611) then return to_sfixed(0.00062073246430788330, 1, -nbits);
    elsif (x=1612) then return to_sfixed(0.00062034739454094293, 1, -nbits);
    elsif (x=1613) then return to_sfixed(0.00061996280223186606, 1, -nbits);
    elsif (x=1614) then return to_sfixed(0.00061957868649318464, 1, -nbits);
    elsif (x=1615) then return to_sfixed(0.00061919504643962852, 1, -nbits);
    elsif (x=1616) then return to_sfixed(0.00061881188118811882, 1, -nbits);
    elsif (x=1617) then return to_sfixed(0.00061842918985776133, 1, -nbits);
    elsif (x=1618) then return to_sfixed(0.00061804697156983925, 1, -nbits);
    elsif (x=1619) then return to_sfixed(0.00061766522544780733, 1, -nbits);
    elsif (x=1620) then return to_sfixed(0.00061728395061728394, 1, -nbits);
    elsif (x=1621) then return to_sfixed(0.00061690314620604567, 1, -nbits);
    elsif (x=1622) then return to_sfixed(0.00061652281134401974, 1, -nbits);
    elsif (x=1623) then return to_sfixed(0.00061614294516327791, 1, -nbits);
    elsif (x=1624) then return to_sfixed(0.00061576354679802956, 1, -nbits);
    elsif (x=1625) then return to_sfixed(0.00061538461538461541, 1, -nbits);
    elsif (x=1626) then return to_sfixed(0.00061500615006150063, 1, -nbits);
    elsif (x=1627) then return to_sfixed(0.00061462814996926854, 1, -nbits);
    elsif (x=1628) then return to_sfixed(0.00061425061425061424, 1, -nbits);
    elsif (x=1629) then return to_sfixed(0.00061387354205033758, 1, -nbits);
    elsif (x=1630) then return to_sfixed(0.00061349693251533746, 1, -nbits);
    elsif (x=1631) then return to_sfixed(0.00061312078479460450, 1, -nbits);
    elsif (x=1632) then return to_sfixed(0.00061274509803921568, 1, -nbits);
    elsif (x=1633) then return to_sfixed(0.00061236987140232701, 1, -nbits);
    elsif (x=1634) then return to_sfixed(0.00061199510403916763, 1, -nbits);
    elsif (x=1635) then return to_sfixed(0.00061162079510703360, 1, -nbits);
    elsif (x=1636) then return to_sfixed(0.00061124694376528117, 1, -nbits);
    elsif (x=1637) then return to_sfixed(0.00061087354917532073, 1, -nbits);
    elsif (x=1638) then return to_sfixed(0.00061050061050061050, 1, -nbits);
    elsif (x=1639) then return to_sfixed(0.00061012812690665037, 1, -nbits);
    elsif (x=1640) then return to_sfixed(0.00060975609756097561, 1, -nbits);
    elsif (x=1641) then return to_sfixed(0.00060938452163315055, 1, -nbits);
    elsif (x=1642) then return to_sfixed(0.00060901339829476245, 1, -nbits);
    elsif (x=1643) then return to_sfixed(0.00060864272671941571, 1, -nbits);
    elsif (x=1644) then return to_sfixed(0.00060827250608272508, 1, -nbits);
    elsif (x=1645) then return to_sfixed(0.00060790273556231007, 1, -nbits);
    elsif (x=1646) then return to_sfixed(0.00060753341433778852, 1, -nbits);
    elsif (x=1647) then return to_sfixed(0.00060716454159077113, 1, -nbits);
    elsif (x=1648) then return to_sfixed(0.00060679611650485432, 1, -nbits);
    elsif (x=1649) then return to_sfixed(0.00060642813826561554, 1, -nbits);
    elsif (x=1650) then return to_sfixed(0.00060606060606060606, 1, -nbits);
    elsif (x=1651) then return to_sfixed(0.00060569351907934583, 1, -nbits);
    elsif (x=1652) then return to_sfixed(0.00060532687651331722, 1, -nbits);
    elsif (x=1653) then return to_sfixed(0.00060496067755595891, 1, -nbits);
    elsif (x=1654) then return to_sfixed(0.00060459492140266019, 1, -nbits);
    elsif (x=1655) then return to_sfixed(0.00060422960725075529, 1, -nbits);
    elsif (x=1656) then return to_sfixed(0.00060386473429951688, 1, -nbits);
    elsif (x=1657) then return to_sfixed(0.00060350030175015089, 1, -nbits);
    elsif (x=1658) then return to_sfixed(0.00060313630880579007, 1, -nbits);
    elsif (x=1659) then return to_sfixed(0.00060277275467148883, 1, -nbits);
    elsif (x=1660) then return to_sfixed(0.00060240963855421692, 1, -nbits);
    elsif (x=1661) then return to_sfixed(0.00060204695966285370, 1, -nbits);
    elsif (x=1662) then return to_sfixed(0.00060168471720818293, 1, -nbits);
    elsif (x=1663) then return to_sfixed(0.00060132291040288638, 1, -nbits);
    elsif (x=1664) then return to_sfixed(0.00060096153846153849, 1, -nbits);
    elsif (x=1665) then return to_sfixed(0.00060060060060060057, 1, -nbits);
    elsif (x=1666) then return to_sfixed(0.00060024009603841532, 1, -nbits);
    elsif (x=1667) then return to_sfixed(0.00059988002399520091, 1, -nbits);
    elsif (x=1668) then return to_sfixed(0.00059952038369304552, 1, -nbits);
    elsif (x=1669) then return to_sfixed(0.00059916117435590175, 1, -nbits);
    elsif (x=1670) then return to_sfixed(0.00059880239520958083, 1, -nbits);
    elsif (x=1671) then return to_sfixed(0.00059844404548174744, 1, -nbits);
    elsif (x=1672) then return to_sfixed(0.00059808612440191385, 1, -nbits);
    elsif (x=1673) then return to_sfixed(0.00059772863120143450, 1, -nbits);
    elsif (x=1674) then return to_sfixed(0.00059737156511350056, 1, -nbits);
    elsif (x=1675) then return to_sfixed(0.00059701492537313433, 1, -nbits);
    elsif (x=1676) then return to_sfixed(0.00059665871121718380, 1, -nbits);
    elsif (x=1677) then return to_sfixed(0.00059630292188431720, 1, -nbits);
    elsif (x=1678) then return to_sfixed(0.00059594755661501785, 1, -nbits);
    elsif (x=1679) then return to_sfixed(0.00059559261465157837, 1, -nbits);
    elsif (x=1680) then return to_sfixed(0.00059523809523809529, 1, -nbits);
    elsif (x=1681) then return to_sfixed(0.00059488399762046404, 1, -nbits);
    elsif (x=1682) then return to_sfixed(0.00059453032104637331, 1, -nbits);
    elsif (x=1683) then return to_sfixed(0.00059417706476530010, 1, -nbits);
    elsif (x=1684) then return to_sfixed(0.00059382422802850359, 1, -nbits);
    elsif (x=1685) then return to_sfixed(0.00059347181008902075, 1, -nbits);
    elsif (x=1686) then return to_sfixed(0.00059311981020166078, 1, -nbits);
    elsif (x=1687) then return to_sfixed(0.00059276822762299936, 1, -nbits);
    elsif (x=1688) then return to_sfixed(0.00059241706161137445, 1, -nbits);
    elsif (x=1689) then return to_sfixed(0.00059206631142687976, 1, -nbits);
    elsif (x=1690) then return to_sfixed(0.00059171597633136095, 1, -nbits);
    elsif (x=1691) then return to_sfixed(0.00059136605558840927, 1, -nbits);
    elsif (x=1692) then return to_sfixed(0.00059101654846335696, 1, -nbits);
    elsif (x=1693) then return to_sfixed(0.00059066745422327229, 1, -nbits);
    elsif (x=1694) then return to_sfixed(0.00059031877213695393, 1, -nbits);
    elsif (x=1695) then return to_sfixed(0.00058997050147492625, 1, -nbits);
    elsif (x=1696) then return to_sfixed(0.00058962264150943394, 1, -nbits);
    elsif (x=1697) then return to_sfixed(0.00058927519151443723, 1, -nbits);
    elsif (x=1698) then return to_sfixed(0.00058892815076560655, 1, -nbits);
    elsif (x=1699) then return to_sfixed(0.00058858151854031780, 1, -nbits);
    elsif (x=1700) then return to_sfixed(0.00058823529411764701, 1, -nbits);
    elsif (x=1701) then return to_sfixed(0.00058788947677836567, 1, -nbits);
    elsif (x=1702) then return to_sfixed(0.00058754406580493535, 1, -nbits);
    elsif (x=1703) then return to_sfixed(0.00058719906048150322, 1, -nbits);
    elsif (x=1704) then return to_sfixed(0.00058685446009389673, 1, -nbits);
    elsif (x=1705) then return to_sfixed(0.00058651026392961877, 1, -nbits);
    elsif (x=1706) then return to_sfixed(0.00058616647127784287, 1, -nbits);
    elsif (x=1707) then return to_sfixed(0.00058582308142940832, 1, -nbits);
    elsif (x=1708) then return to_sfixed(0.00058548009367681499, 1, -nbits);
    elsif (x=1709) then return to_sfixed(0.00058513750731421885, 1, -nbits);
    elsif (x=1710) then return to_sfixed(0.00058479532163742691, 1, -nbits);
    elsif (x=1711) then return to_sfixed(0.00058445353594389242, 1, -nbits);
    elsif (x=1712) then return to_sfixed(0.00058411214953271024, 1, -nbits);
    elsif (x=1713) then return to_sfixed(0.00058377116170461180, 1, -nbits);
    elsif (x=1714) then return to_sfixed(0.00058343057176196028, 1, -nbits);
    elsif (x=1715) then return to_sfixed(0.00058309037900874635, 1, -nbits);
    elsif (x=1716) then return to_sfixed(0.00058275058275058275, 1, -nbits);
    elsif (x=1717) then return to_sfixed(0.00058241118229470008, 1, -nbits);
    elsif (x=1718) then return to_sfixed(0.00058207217694994178, 1, -nbits);
    elsif (x=1719) then return to_sfixed(0.00058173356602675972, 1, -nbits);
    elsif (x=1720) then return to_sfixed(0.00058139534883720929, 1, -nbits);
    elsif (x=1721) then return to_sfixed(0.00058105752469494478, 1, -nbits);
    elsif (x=1722) then return to_sfixed(0.00058072009291521487, 1, -nbits);
    elsif (x=1723) then return to_sfixed(0.00058038305281485781, 1, -nbits);
    elsif (x=1724) then return to_sfixed(0.00058004640371229696, 1, -nbits);
    elsif (x=1725) then return to_sfixed(0.00057971014492753622, 1, -nbits);
    elsif (x=1726) then return to_sfixed(0.00057937427578215526, 1, -nbits);
    elsif (x=1727) then return to_sfixed(0.00057903879559930511, 1, -nbits);
    elsif (x=1728) then return to_sfixed(0.00057870370370370367, 1, -nbits);
    elsif (x=1729) then return to_sfixed(0.00057836899942163096, 1, -nbits);
    elsif (x=1730) then return to_sfixed(0.00057803468208092489, 1, -nbits);
    elsif (x=1731) then return to_sfixed(0.00057770075101097628, 1, -nbits);
    elsif (x=1732) then return to_sfixed(0.00057736720554272516, 1, -nbits);
    elsif (x=1733) then return to_sfixed(0.00057703404500865547, 1, -nbits);
    elsif (x=1734) then return to_sfixed(0.00057670126874279125, 1, -nbits);
    elsif (x=1735) then return to_sfixed(0.00057636887608069167, 1, -nbits);
    elsif (x=1736) then return to_sfixed(0.00057603686635944700, 1, -nbits);
    elsif (x=1737) then return to_sfixed(0.00057570523891767420, 1, -nbits);
    elsif (x=1738) then return to_sfixed(0.00057537399309551208, 1, -nbits);
    elsif (x=1739) then return to_sfixed(0.00057504312823461760, 1, -nbits);
    elsif (x=1740) then return to_sfixed(0.00057471264367816091, 1, -nbits);
    elsif (x=1741) then return to_sfixed(0.00057438253877082138, 1, -nbits);
    elsif (x=1742) then return to_sfixed(0.00057405281285878302, 1, -nbits);
    elsif (x=1743) then return to_sfixed(0.00057372346528973030, 1, -nbits);
    elsif (x=1744) then return to_sfixed(0.00057339449541284407, 1, -nbits);
    elsif (x=1745) then return to_sfixed(0.00057306590257879652, 1, -nbits);
    elsif (x=1746) then return to_sfixed(0.00057273768613974802, 1, -nbits);
    elsif (x=1747) then return to_sfixed(0.00057240984544934168, 1, -nbits);
    elsif (x=1748) then return to_sfixed(0.00057208237986270023, 1, -nbits);
    elsif (x=1749) then return to_sfixed(0.00057175528873642080, 1, -nbits);
    elsif (x=1750) then return to_sfixed(0.00057142857142857147, 1, -nbits);
    elsif (x=1751) then return to_sfixed(0.00057110222729868647, 1, -nbits);
    elsif (x=1752) then return to_sfixed(0.00057077625570776253, 1, -nbits);
    elsif (x=1753) then return to_sfixed(0.00057045065601825438, 1, -nbits);
    elsif (x=1754) then return to_sfixed(0.00057012542759407071, 1, -nbits);
    elsif (x=1755) then return to_sfixed(0.00056980056980056976, 1, -nbits);
    elsif (x=1756) then return to_sfixed(0.00056947608200455578, 1, -nbits);
    elsif (x=1757) then return to_sfixed(0.00056915196357427435, 1, -nbits);
    elsif (x=1758) then return to_sfixed(0.00056882821387940839, 1, -nbits);
    elsif (x=1759) then return to_sfixed(0.00056850483229107444, 1, -nbits);
    elsif (x=1760) then return to_sfixed(0.00056818181818181815, 1, -nbits);
    elsif (x=1761) then return to_sfixed(0.00056785917092561046, 1, -nbits);
    elsif (x=1762) then return to_sfixed(0.00056753688989784334, 1, -nbits);
    elsif (x=1763) then return to_sfixed(0.00056721497447532619, 1, -nbits);
    elsif (x=1764) then return to_sfixed(0.00056689342403628119, 1, -nbits);
    elsif (x=1765) then return to_sfixed(0.00056657223796033991, 1, -nbits);
    elsif (x=1766) then return to_sfixed(0.00056625141562853911, 1, -nbits);
    elsif (x=1767) then return to_sfixed(0.00056593095642331638, 1, -nbits);
    elsif (x=1768) then return to_sfixed(0.00056561085972850684, 1, -nbits);
    elsif (x=1769) then return to_sfixed(0.00056529112492933857, 1, -nbits);
    elsif (x=1770) then return to_sfixed(0.00056497175141242940, 1, -nbits);
    elsif (x=1771) then return to_sfixed(0.00056465273856578201, 1, -nbits);
    elsif (x=1772) then return to_sfixed(0.00056433408577878099, 1, -nbits);
    elsif (x=1773) then return to_sfixed(0.00056401579244218843, 1, -nbits);
    elsif (x=1774) then return to_sfixed(0.00056369785794813977, 1, -nbits);
    elsif (x=1775) then return to_sfixed(0.00056338028169014088, 1, -nbits);
    elsif (x=1776) then return to_sfixed(0.00056306306306306306, 1, -nbits);
    elsif (x=1777) then return to_sfixed(0.00056274620146314015, 1, -nbits);
    elsif (x=1778) then return to_sfixed(0.00056242969628796406, 1, -nbits);
    elsif (x=1779) then return to_sfixed(0.00056211354693648118, 1, -nbits);
    elsif (x=1780) then return to_sfixed(0.00056179775280898881, 1, -nbits);
    elsif (x=1781) then return to_sfixed(0.00056148231330713087, 1, -nbits);
    elsif (x=1782) then return to_sfixed(0.00056116722783389455, 1, -nbits);
    elsif (x=1783) then return to_sfixed(0.00056085249579360629, 1, -nbits);
    elsif (x=1784) then return to_sfixed(0.00056053811659192824, 1, -nbits);
    elsif (x=1785) then return to_sfixed(0.00056022408963585430, 1, -nbits);
    elsif (x=1786) then return to_sfixed(0.00055991041433370661, 1, -nbits);
    elsif (x=1787) then return to_sfixed(0.00055959709009513155, 1, -nbits);
    elsif (x=1788) then return to_sfixed(0.00055928411633109618, 1, -nbits);
    elsif (x=1789) then return to_sfixed(0.00055897149245388487, 1, -nbits);
    elsif (x=1790) then return to_sfixed(0.00055865921787709492, 1, -nbits);
    elsif (x=1791) then return to_sfixed(0.00055834729201563373, 1, -nbits);
    elsif (x=1792) then return to_sfixed(0.00055803571428571425, 1, -nbits);
    elsif (x=1793) then return to_sfixed(0.00055772448410485224, 1, -nbits);
    elsif (x=1794) then return to_sfixed(0.00055741360089186175, 1, -nbits);
    elsif (x=1795) then return to_sfixed(0.00055710306406685239, 1, -nbits);
    elsif (x=1796) then return to_sfixed(0.00055679287305122492, 1, -nbits);
    elsif (x=1797) then return to_sfixed(0.00055648302726766835, 1, -nbits);
    elsif (x=1798) then return to_sfixed(0.00055617352614015572, 1, -nbits);
    elsif (x=1799) then return to_sfixed(0.00055586436909394106, 1, -nbits);
    elsif (x=1800) then return to_sfixed(0.00055555555555555556, 1, -nbits);
    elsif (x=1801) then return to_sfixed(0.00055524708495280405, 1, -nbits);
    elsif (x=1802) then return to_sfixed(0.00055493895671476139, 1, -nbits);
    elsif (x=1803) then return to_sfixed(0.00055463117027176932, 1, -nbits);
    elsif (x=1804) then return to_sfixed(0.00055432372505543237, 1, -nbits);
    elsif (x=1805) then return to_sfixed(0.00055401662049861500, 1, -nbits);
    elsif (x=1806) then return to_sfixed(0.00055370985603543741, 1, -nbits);
    elsif (x=1807) then return to_sfixed(0.00055340343110127279, 1, -nbits);
    elsif (x=1808) then return to_sfixed(0.00055309734513274336, 1, -nbits);
    elsif (x=1809) then return to_sfixed(0.00055279159756771695, 1, -nbits);
    elsif (x=1810) then return to_sfixed(0.00055248618784530391, 1, -nbits);
    elsif (x=1811) then return to_sfixed(0.00055218111540585317, 1, -nbits);
    elsif (x=1812) then return to_sfixed(0.00055187637969094923, 1, -nbits);
    elsif (x=1813) then return to_sfixed(0.00055157198014340876, 1, -nbits);
    elsif (x=1814) then return to_sfixed(0.00055126791620727675, 1, -nbits);
    elsif (x=1815) then return to_sfixed(0.00055096418732782364, 1, -nbits);
    elsif (x=1816) then return to_sfixed(0.00055066079295154190, 1, -nbits);
    elsif (x=1817) then return to_sfixed(0.00055035773252614197, 1, -nbits);
    elsif (x=1818) then return to_sfixed(0.00055005500550055003, 1, -nbits);
    elsif (x=1819) then return to_sfixed(0.00054975261132490382, 1, -nbits);
    elsif (x=1820) then return to_sfixed(0.00054945054945054945, 1, -nbits);
    elsif (x=1821) then return to_sfixed(0.00054914881933003845, 1, -nbits);
    elsif (x=1822) then return to_sfixed(0.00054884742041712406, 1, -nbits);
    elsif (x=1823) then return to_sfixed(0.00054854635216675812, 1, -nbits);
    elsif (x=1824) then return to_sfixed(0.00054824561403508769, 1, -nbits);
    elsif (x=1825) then return to_sfixed(0.00054794520547945202, 1, -nbits);
    elsif (x=1826) then return to_sfixed(0.00054764512595837896, 1, -nbits);
    elsif (x=1827) then return to_sfixed(0.00054734537493158185, 1, -nbits);
    elsif (x=1828) then return to_sfixed(0.00054704595185995622, 1, -nbits);
    elsif (x=1829) then return to_sfixed(0.00054674685620557679, 1, -nbits);
    elsif (x=1830) then return to_sfixed(0.00054644808743169399, 1, -nbits);
    elsif (x=1831) then return to_sfixed(0.00054614964500273070, 1, -nbits);
    elsif (x=1832) then return to_sfixed(0.00054585152838427945, 1, -nbits);
    elsif (x=1833) then return to_sfixed(0.00054555373704309870, 1, -nbits);
    elsif (x=1834) then return to_sfixed(0.00054525627044711017, 1, -nbits);
    elsif (x=1835) then return to_sfixed(0.00054495912806539512, 1, -nbits);
    elsif (x=1836) then return to_sfixed(0.00054466230936819177, 1, -nbits);
    elsif (x=1837) then return to_sfixed(0.00054436581382689172, 1, -nbits);
    elsif (x=1838) then return to_sfixed(0.00054406964091403701, 1, -nbits);
    elsif (x=1839) then return to_sfixed(0.00054377379010331697, 1, -nbits);
    elsif (x=1840) then return to_sfixed(0.00054347826086956522, 1, -nbits);
    elsif (x=1841) then return to_sfixed(0.00054318305268875606, 1, -nbits);
    elsif (x=1842) then return to_sfixed(0.00054288816503800220, 1, -nbits);
    elsif (x=1843) then return to_sfixed(0.00054259359739555074, 1, -nbits);
    elsif (x=1844) then return to_sfixed(0.00054229934924078093, 1, -nbits);
    elsif (x=1845) then return to_sfixed(0.00054200542005420054, 1, -nbits);
    elsif (x=1846) then return to_sfixed(0.00054171180931744309, 1, -nbits);
    elsif (x=1847) then return to_sfixed(0.00054141851651326478, 1, -nbits);
    elsif (x=1848) then return to_sfixed(0.00054112554112554113, 1, -nbits);
    elsif (x=1849) then return to_sfixed(0.00054083288263926451, 1, -nbits);
    elsif (x=1850) then return to_sfixed(0.00054054054054054055, 1, -nbits);
    elsif (x=1851) then return to_sfixed(0.00054024851431658564, 1, -nbits);
    elsif (x=1852) then return to_sfixed(0.00053995680345572358, 1, -nbits);
    elsif (x=1853) then return to_sfixed(0.00053966540744738263, 1, -nbits);
    elsif (x=1854) then return to_sfixed(0.00053937432578209273, 1, -nbits);
    elsif (x=1855) then return to_sfixed(0.00053908355795148253, 1, -nbits);
    elsif (x=1856) then return to_sfixed(0.00053879310344827585, 1, -nbits);
    elsif (x=1857) then return to_sfixed(0.00053850296176628971, 1, -nbits);
    elsif (x=1858) then return to_sfixed(0.00053821313240043052, 1, -nbits);
    elsif (x=1859) then return to_sfixed(0.00053792361484669173, 1, -nbits);
    elsif (x=1860) then return to_sfixed(0.00053763440860215054, 1, -nbits);
    elsif (x=1861) then return to_sfixed(0.00053734551316496511, 1, -nbits);
    elsif (x=1862) then return to_sfixed(0.00053705692803437163, 1, -nbits);
    elsif (x=1863) then return to_sfixed(0.00053676865271068169, 1, -nbits);
    elsif (x=1864) then return to_sfixed(0.00053648068669527897, 1, -nbits);
    elsif (x=1865) then return to_sfixed(0.00053619302949061668, 1, -nbits);
    elsif (x=1866) then return to_sfixed(0.00053590568060021436, 1, -nbits);
    elsif (x=1867) then return to_sfixed(0.00053561863952865559, 1, -nbits);
    elsif (x=1868) then return to_sfixed(0.00053533190578158461, 1, -nbits);
    elsif (x=1869) then return to_sfixed(0.00053504547886570354, 1, -nbits);
    elsif (x=1870) then return to_sfixed(0.00053475935828877007, 1, -nbits);
    elsif (x=1871) then return to_sfixed(0.00053447354355959376, 1, -nbits);
    elsif (x=1872) then return to_sfixed(0.00053418803418803424, 1, -nbits);
    elsif (x=1873) then return to_sfixed(0.00053390282968499730, 1, -nbits);
    elsif (x=1874) then return to_sfixed(0.00053361792956243333, 1, -nbits);
    elsif (x=1875) then return to_sfixed(0.00053333333333333336, 1, -nbits);
    elsif (x=1876) then return to_sfixed(0.00053304904051172707, 1, -nbits);
    elsif (x=1877) then return to_sfixed(0.00053276505061267978, 1, -nbits);
    elsif (x=1878) then return to_sfixed(0.00053248136315228972, 1, -nbits);
    elsif (x=1879) then return to_sfixed(0.00053219797764768491, 1, -nbits);
    elsif (x=1880) then return to_sfixed(0.00053191489361702129, 1, -nbits);
    elsif (x=1881) then return to_sfixed(0.00053163211057947904, 1, -nbits);
    elsif (x=1882) then return to_sfixed(0.00053134962805526033, 1, -nbits);
    elsif (x=1883) then return to_sfixed(0.00053106744556558679, 1, -nbits);
    elsif (x=1884) then return to_sfixed(0.00053078556263269638, 1, -nbits);
    elsif (x=1885) then return to_sfixed(0.00053050397877984080, 1, -nbits);
    elsif (x=1886) then return to_sfixed(0.00053022269353128319, 1, -nbits);
    elsif (x=1887) then return to_sfixed(0.00052994170641229468, 1, -nbits);
    elsif (x=1888) then return to_sfixed(0.00052966101694915254, 1, -nbits);
    elsif (x=1889) then return to_sfixed(0.00052938062466913714, 1, -nbits);
    elsif (x=1890) then return to_sfixed(0.00052910052910052914, 1, -nbits);
    elsif (x=1891) then return to_sfixed(0.00052882072977260709, 1, -nbits);
    elsif (x=1892) then return to_sfixed(0.00052854122621564484, 1, -nbits);
    elsif (x=1893) then return to_sfixed(0.00052826201796090863, 1, -nbits);
    elsif (x=1894) then return to_sfixed(0.00052798310454065466, 1, -nbits);
    elsif (x=1895) then return to_sfixed(0.00052770448548812663, 1, -nbits);
    elsif (x=1896) then return to_sfixed(0.00052742616033755270, 1, -nbits);
    elsif (x=1897) then return to_sfixed(0.00052714812862414342, 1, -nbits);
    elsif (x=1898) then return to_sfixed(0.00052687038988408848, 1, -nbits);
    elsif (x=1899) then return to_sfixed(0.00052659294365455498, 1, -nbits);
    elsif (x=1900) then return to_sfixed(0.00052631578947368420, 1, -nbits);
    elsif (x=1901) then return to_sfixed(0.00052603892688058915, 1, -nbits);
    elsif (x=1902) then return to_sfixed(0.00052576235541535224, 1, -nbits);
    elsif (x=1903) then return to_sfixed(0.00052548607461902258, 1, -nbits);
    elsif (x=1904) then return to_sfixed(0.00052521008403361342, 1, -nbits);
    elsif (x=1905) then return to_sfixed(0.00052493438320209973, 1, -nbits);
    elsif (x=1906) then return to_sfixed(0.00052465897166841555, 1, -nbits);
    elsif (x=1907) then return to_sfixed(0.00052438384897745150, 1, -nbits);
    elsif (x=1908) then return to_sfixed(0.00052410901467505244, 1, -nbits);
    elsif (x=1909) then return to_sfixed(0.00052383446830801469, 1, -nbits);
    elsif (x=1910) then return to_sfixed(0.00052356020942408382, 1, -nbits);
    elsif (x=1911) then return to_sfixed(0.00052328623757195189, 1, -nbits);
    elsif (x=1912) then return to_sfixed(0.00052301255230125519, 1, -nbits);
    elsif (x=1913) then return to_sfixed(0.00052273915316257186, 1, -nbits);
    elsif (x=1914) then return to_sfixed(0.00052246603970741907, 1, -nbits);
    elsif (x=1915) then return to_sfixed(0.00052219321148825064, 1, -nbits);
    elsif (x=1916) then return to_sfixed(0.00052192066805845506, 1, -nbits);
    elsif (x=1917) then return to_sfixed(0.00052164840897235261, 1, -nbits);
    elsif (x=1918) then return to_sfixed(0.00052137643378519292, 1, -nbits);
    elsif (x=1919) then return to_sfixed(0.00052110474205315264, 1, -nbits);
    elsif (x=1920) then return to_sfixed(0.00052083333333333333, 1, -nbits);
    elsif (x=1921) then return to_sfixed(0.00052056220718375845, 1, -nbits);
    elsif (x=1922) then return to_sfixed(0.00052029136316337154, 1, -nbits);
    elsif (x=1923) then return to_sfixed(0.00052002080083203334, 1, -nbits);
    elsif (x=1924) then return to_sfixed(0.00051975051975051978, 1, -nbits);
    elsif (x=1925) then return to_sfixed(0.00051948051948051948, 1, -nbits);
    elsif (x=1926) then return to_sfixed(0.00051921079958463135, 1, -nbits);
    elsif (x=1927) then return to_sfixed(0.00051894135962636220, 1, -nbits);
    elsif (x=1928) then return to_sfixed(0.00051867219917012448, 1, -nbits);
    elsif (x=1929) then return to_sfixed(0.00051840331778123380, 1, -nbits);
    elsif (x=1930) then return to_sfixed(0.00051813471502590671, 1, -nbits);
    elsif (x=1931) then return to_sfixed(0.00051786639047125837, 1, -nbits);
    elsif (x=1932) then return to_sfixed(0.00051759834368530024, 1, -nbits);
    elsif (x=1933) then return to_sfixed(0.00051733057423693739, 1, -nbits);
    elsif (x=1934) then return to_sfixed(0.00051706308169596695, 1, -nbits);
    elsif (x=1935) then return to_sfixed(0.00051679586563307489, 1, -nbits);
    elsif (x=1936) then return to_sfixed(0.00051652892561983473, 1, -nbits);
    elsif (x=1937) then return to_sfixed(0.00051626226122870422, 1, -nbits);
    elsif (x=1938) then return to_sfixed(0.00051599587203302369, 1, -nbits);
    elsif (x=1939) then return to_sfixed(0.00051572975760701394, 1, -nbits);
    elsif (x=1940) then return to_sfixed(0.00051546391752577321, 1, -nbits);
    elsif (x=1941) then return to_sfixed(0.00051519835136527566, 1, -nbits);
    elsif (x=1942) then return to_sfixed(0.00051493305870236867, 1, -nbits);
    elsif (x=1943) then return to_sfixed(0.00051466803911477102, 1, -nbits);
    elsif (x=1944) then return to_sfixed(0.00051440329218107000, 1, -nbits);
    elsif (x=1945) then return to_sfixed(0.00051413881748071976, 1, -nbits);
    elsif (x=1946) then return to_sfixed(0.00051387461459403907, 1, -nbits);
    elsif (x=1947) then return to_sfixed(0.00051361068310220854, 1, -nbits);
    elsif (x=1948) then return to_sfixed(0.00051334702258726901, 1, -nbits);
    elsif (x=1949) then return to_sfixed(0.00051308363263211901, 1, -nbits);
    elsif (x=1950) then return to_sfixed(0.00051282051282051282, 1, -nbits);
    elsif (x=1951) then return to_sfixed(0.00051255766273705791, 1, -nbits);
    elsif (x=1952) then return to_sfixed(0.00051229508196721314, 1, -nbits);
    elsif (x=1953) then return to_sfixed(0.00051203277009728623, 1, -nbits);
    elsif (x=1954) then return to_sfixed(0.00051177072671443195, 1, -nbits);
    elsif (x=1955) then return to_sfixed(0.00051150895140664957, 1, -nbits);
    elsif (x=1956) then return to_sfixed(0.00051124744376278123, 1, -nbits);
    elsif (x=1957) then return to_sfixed(0.00051098620337250899, 1, -nbits);
    elsif (x=1958) then return to_sfixed(0.00051072522982635344, 1, -nbits);
    elsif (x=1959) then return to_sfixed(0.00051046452271567128, 1, -nbits);
    elsif (x=1960) then return to_sfixed(0.00051020408163265311, 1, -nbits);
    elsif (x=1961) then return to_sfixed(0.00050994390617032130, 1, -nbits);
    elsif (x=1962) then return to_sfixed(0.00050968399592252807, 1, -nbits);
    elsif (x=1963) then return to_sfixed(0.00050942435048395313, 1, -nbits);
    elsif (x=1964) then return to_sfixed(0.00050916496945010179, 1, -nbits);
    elsif (x=1965) then return to_sfixed(0.00050890585241730279, 1, -nbits);
    elsif (x=1966) then return to_sfixed(0.00050864699898270599, 1, -nbits);
    elsif (x=1967) then return to_sfixed(0.00050838840874428064, 1, -nbits);
    elsif (x=1968) then return to_sfixed(0.00050813008130081306, 1, -nbits);
    elsif (x=1969) then return to_sfixed(0.00050787201625190448, 1, -nbits);
    elsif (x=1970) then return to_sfixed(0.00050761421319796957, 1, -nbits);
    elsif (x=1971) then return to_sfixed(0.00050735667174023336, 1, -nbits);
    elsif (x=1972) then return to_sfixed(0.00050709939148073022, 1, -nbits);
    elsif (x=1973) then return to_sfixed(0.00050684237202230106, 1, -nbits);
    elsif (x=1974) then return to_sfixed(0.00050658561296859173, 1, -nbits);
    elsif (x=1975) then return to_sfixed(0.00050632911392405066, 1, -nbits);
    elsif (x=1976) then return to_sfixed(0.00050607287449392713, 1, -nbits);
    elsif (x=1977) then return to_sfixed(0.00050581689428426911, 1, -nbits);
    elsif (x=1978) then return to_sfixed(0.00050556117290192115, 1, -nbits);
    elsif (x=1979) then return to_sfixed(0.00050530570995452253, 1, -nbits);
    elsif (x=1980) then return to_sfixed(0.00050505050505050505, 1, -nbits);
    elsif (x=1981) then return to_sfixed(0.00050479555779909136, 1, -nbits);
    elsif (x=1982) then return to_sfixed(0.00050454086781029264, 1, -nbits);
    elsif (x=1983) then return to_sfixed(0.00050428643469490675, 1, -nbits);
    elsif (x=1984) then return to_sfixed(0.00050403225806451612, 1, -nbits);
    elsif (x=1985) then return to_sfixed(0.00050377833753148613, 1, -nbits);
    elsif (x=1986) then return to_sfixed(0.00050352467270896274, 1, -nbits);
    elsif (x=1987) then return to_sfixed(0.00050327126321087065, 1, -nbits);
    elsif (x=1988) then return to_sfixed(0.00050301810865191151, 1, -nbits);
    elsif (x=1989) then return to_sfixed(0.00050276520864756154, 1, -nbits);
    elsif (x=1990) then return to_sfixed(0.00050251256281407040, 1, -nbits);
    elsif (x=1991) then return to_sfixed(0.00050226017076845811, 1, -nbits);
    elsif (x=1992) then return to_sfixed(0.00050200803212851401, 1, -nbits);
    elsif (x=1993) then return to_sfixed(0.00050175614651279475, 1, -nbits);
    elsif (x=1994) then return to_sfixed(0.00050150451354062187, 1, -nbits);
    elsif (x=1995) then return to_sfixed(0.00050125313283208019, 1, -nbits);
    elsif (x=1996) then return to_sfixed(0.00050100200400801599, 1, -nbits);
    elsif (x=1997) then return to_sfixed(0.00050075112669003500, 1, -nbits);
    elsif (x=1998) then return to_sfixed(0.00050050050050050050, 1, -nbits);
    elsif (x=1999) then return to_sfixed(0.00050025012506253123, 1, -nbits);
    elsif (x=2000) then return to_sfixed(0.00050000000000000001, 1, -nbits);
    elsif (x=2001) then return to_sfixed(0.00049975012493753122, 1, -nbits);
    elsif (x=2002) then return to_sfixed(0.00049950049950049950, 1, -nbits);
    elsif (x=2003) then return to_sfixed(0.00049925112331502750, 1, -nbits);
    elsif (x=2004) then return to_sfixed(0.00049900199600798399, 1, -nbits);
    elsif (x=2005) then return to_sfixed(0.00049875311720698251, 1, -nbits);
    elsif (x=2006) then return to_sfixed(0.00049850448654037882, 1, -nbits);
    elsif (x=2007) then return to_sfixed(0.00049825610363726954, 1, -nbits);
    elsif (x=2008) then return to_sfixed(0.00049800796812749003, 1, -nbits);
    elsif (x=2009) then return to_sfixed(0.00049776007964161273, 1, -nbits);
    elsif (x=2010) then return to_sfixed(0.00049751243781094524, 1, -nbits);
    elsif (x=2011) then return to_sfixed(0.00049726504226752855, 1, -nbits);
    elsif (x=2012) then return to_sfixed(0.00049701789264413514, 1, -nbits);
    elsif (x=2013) then return to_sfixed(0.00049677098857426726, 1, -nbits);
    elsif (x=2014) then return to_sfixed(0.00049652432969215490, 1, -nbits);
    elsif (x=2015) then return to_sfixed(0.00049627791563275434, 1, -nbits);
    elsif (x=2016) then return to_sfixed(0.00049603174603174600, 1, -nbits);
    elsif (x=2017) then return to_sfixed(0.00049578582052553293, 1, -nbits);
    elsif (x=2018) then return to_sfixed(0.00049554013875123884, 1, -nbits);
    elsif (x=2019) then return to_sfixed(0.00049529470034670627, 1, -nbits);
    elsif (x=2020) then return to_sfixed(0.00049504950495049506, 1, -nbits);
    elsif (x=2021) then return to_sfixed(0.00049480455220188031, 1, -nbits);
    elsif (x=2022) then return to_sfixed(0.00049455984174085062, 1, -nbits);
    elsif (x=2023) then return to_sfixed(0.00049431537320810673, 1, -nbits);
    elsif (x=2024) then return to_sfixed(0.00049407114624505926, 1, -nbits);
    elsif (x=2025) then return to_sfixed(0.00049382716049382717, 1, -nbits);
    elsif (x=2026) then return to_sfixed(0.00049358341559723590, 1, -nbits);
    elsif (x=2027) then return to_sfixed(0.00049333991119881603, 1, -nbits);
    elsif (x=2028) then return to_sfixed(0.00049309664694280081, 1, -nbits);
    elsif (x=2029) then return to_sfixed(0.00049285362247412522, 1, -nbits);
    elsif (x=2030) then return to_sfixed(0.00049261083743842361, 1, -nbits);
    elsif (x=2031) then return to_sfixed(0.00049236829148202859, 1, -nbits);
    elsif (x=2032) then return to_sfixed(0.00049212598425196850, 1, -nbits);
    elsif (x=2033) then return to_sfixed(0.00049188391539596653, 1, -nbits);
    elsif (x=2034) then return to_sfixed(0.00049164208456243857, 1, -nbits);
    elsif (x=2035) then return to_sfixed(0.00049140049140049139, 1, -nbits);
    elsif (x=2036) then return to_sfixed(0.00049115913555992138, 1, -nbits);
    elsif (x=2037) then return to_sfixed(0.00049091801669121256, 1, -nbits);
    elsif (x=2038) then return to_sfixed(0.00049067713444553480, 1, -nbits);
    elsif (x=2039) then return to_sfixed(0.00049043648847474255, 1, -nbits);
    elsif (x=2040) then return to_sfixed(0.00049019607843137254, 1, -nbits);
    elsif (x=2041) then return to_sfixed(0.00048995590396864281, 1, -nbits);
    elsif (x=2042) then return to_sfixed(0.00048971596474045055, 1, -nbits);
    elsif (x=2043) then return to_sfixed(0.00048947626040137058, 1, -nbits);
    elsif (x=2044) then return to_sfixed(0.00048923679060665359, 1, -nbits);
    elsif (x=2045) then return to_sfixed(0.00048899755501222489, 1, -nbits);
    elsif (x=2046) then return to_sfixed(0.00048875855327468231, 1, -nbits);
    elsif (x=2047) then return to_sfixed(0.00048851978505129456, 1, -nbits);
    end if;
  end;


  function reciprocal6 (x : integer; nbits : integer) return sfixed is
  begin
    if (x<1 or x> 6) then
      assert false report "invalid reciprocal6 lookup x=" & integer'image(x) severity warning;
      return to_sfixed(0, 1, -nbits);
    elsif (x=1) then return to_sfixed(1.000000000000, 1, -nbits);
    elsif (x=2) then return to_sfixed(0.500000000000, 1, -nbits);
    elsif (x=3) then return to_sfixed(0.333333333333, 1, -nbits);
    elsif (x=4) then return to_sfixed(0.250000000000, 1, -nbits);
    elsif (x=5) then return to_sfixed(0.200000000000, 1, -nbits);
    elsif (x=6) then return to_sfixed(0.166666666667, 1, -nbits);
    end if;
  end;

end package body reciprocal_pkg;
