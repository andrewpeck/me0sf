library ieee;
use ieee.fixed_pkg.all;

package reciprocal_pkg is
  function reciprocal (x : integer) return sfixed;
end package reciprocal_pkg;

package body reciprocal_pkg is
  --------------------------------------------------------------------------------
  -- functions
  --------------------------------------------------------------------------------


  function reciprocal (x : integer) return sfixed is
  begin
    if (x<1 or x> 630) then
      assert false report "invalid reciprocal lookup x=" & integer'image(x) severity error;
      return to_sfixed(0, 11, -12);
    elsif (x=1) then return to_sfixed(1.000000000000, 11, -12);
    elsif (x=2) then return to_sfixed(0.500000000000, 11, -12);
    elsif (x=3) then return to_sfixed(0.333333333333, 11, -12);
    elsif (x=4) then return to_sfixed(0.250000000000, 11, -12);
    elsif (x=5) then return to_sfixed(0.200000000000, 11, -12);
    elsif (x=6) then return to_sfixed(0.166666666667, 11, -12);
    elsif (x=7) then return to_sfixed(0.142857142857, 11, -12);
    elsif (x=8) then return to_sfixed(0.125000000000, 11, -12);
    elsif (x=9) then return to_sfixed(0.111111111111, 11, -12);
    elsif (x=10) then return to_sfixed(0.100000000000, 11, -12);
    elsif (x=11) then return to_sfixed(0.090909090909, 11, -12);
    elsif (x=12) then return to_sfixed(0.083333333333, 11, -12);
    elsif (x=13) then return to_sfixed(0.076923076923, 11, -12);
    elsif (x=14) then return to_sfixed(0.071428571429, 11, -12);
    elsif (x=15) then return to_sfixed(0.066666666667, 11, -12);
    elsif (x=16) then return to_sfixed(0.062500000000, 11, -12);
    elsif (x=17) then return to_sfixed(0.058823529412, 11, -12);
    elsif (x=18) then return to_sfixed(0.055555555556, 11, -12);
    elsif (x=19) then return to_sfixed(0.052631578947, 11, -12);
    elsif (x=20) then return to_sfixed(0.050000000000, 11, -12);
    elsif (x=21) then return to_sfixed(0.047619047619, 11, -12);
    elsif (x=22) then return to_sfixed(0.045454545455, 11, -12);
    elsif (x=23) then return to_sfixed(0.043478260870, 11, -12);
    elsif (x=24) then return to_sfixed(0.041666666667, 11, -12);
    elsif (x=25) then return to_sfixed(0.040000000000, 11, -12);
    elsif (x=26) then return to_sfixed(0.038461538462, 11, -12);
    elsif (x=27) then return to_sfixed(0.037037037037, 11, -12);
    elsif (x=28) then return to_sfixed(0.035714285714, 11, -12);
    elsif (x=29) then return to_sfixed(0.034482758621, 11, -12);
    elsif (x=30) then return to_sfixed(0.033333333333, 11, -12);
    elsif (x=31) then return to_sfixed(0.032258064516, 11, -12);
    elsif (x=32) then return to_sfixed(0.031250000000, 11, -12);
    elsif (x=33) then return to_sfixed(0.030303030303, 11, -12);
    elsif (x=34) then return to_sfixed(0.029411764706, 11, -12);
    elsif (x=35) then return to_sfixed(0.028571428571, 11, -12);
    elsif (x=36) then return to_sfixed(0.027777777778, 11, -12);
    elsif (x=37) then return to_sfixed(0.027027027027, 11, -12);
    elsif (x=38) then return to_sfixed(0.026315789474, 11, -12);
    elsif (x=39) then return to_sfixed(0.025641025641, 11, -12);
    elsif (x=40) then return to_sfixed(0.025000000000, 11, -12);
    elsif (x=41) then return to_sfixed(0.024390243902, 11, -12);
    elsif (x=42) then return to_sfixed(0.023809523810, 11, -12);
    elsif (x=43) then return to_sfixed(0.023255813953, 11, -12);
    elsif (x=44) then return to_sfixed(0.022727272727, 11, -12);
    elsif (x=45) then return to_sfixed(0.022222222222, 11, -12);
    elsif (x=46) then return to_sfixed(0.021739130435, 11, -12);
    elsif (x=47) then return to_sfixed(0.021276595745, 11, -12);
    elsif (x=48) then return to_sfixed(0.020833333333, 11, -12);
    elsif (x=49) then return to_sfixed(0.020408163265, 11, -12);
    elsif (x=50) then return to_sfixed(0.020000000000, 11, -12);
    elsif (x=51) then return to_sfixed(0.019607843137, 11, -12);
    elsif (x=52) then return to_sfixed(0.019230769231, 11, -12);
    elsif (x=53) then return to_sfixed(0.018867924528, 11, -12);
    elsif (x=54) then return to_sfixed(0.018518518519, 11, -12);
    elsif (x=55) then return to_sfixed(0.018181818182, 11, -12);
    elsif (x=56) then return to_sfixed(0.017857142857, 11, -12);
    elsif (x=57) then return to_sfixed(0.017543859649, 11, -12);
    elsif (x=58) then return to_sfixed(0.017241379310, 11, -12);
    elsif (x=59) then return to_sfixed(0.016949152542, 11, -12);
    elsif (x=60) then return to_sfixed(0.016666666667, 11, -12);
    elsif (x=61) then return to_sfixed(0.016393442623, 11, -12);
    elsif (x=62) then return to_sfixed(0.016129032258, 11, -12);
    elsif (x=63) then return to_sfixed(0.015873015873, 11, -12);
    elsif (x=64) then return to_sfixed(0.015625000000, 11, -12);
    elsif (x=65) then return to_sfixed(0.015384615385, 11, -12);
    elsif (x=66) then return to_sfixed(0.015151515152, 11, -12);
    elsif (x=67) then return to_sfixed(0.014925373134, 11, -12);
    elsif (x=68) then return to_sfixed(0.014705882353, 11, -12);
    elsif (x=69) then return to_sfixed(0.014492753623, 11, -12);
    elsif (x=70) then return to_sfixed(0.014285714286, 11, -12);
    elsif (x=71) then return to_sfixed(0.014084507042, 11, -12);
    elsif (x=72) then return to_sfixed(0.013888888889, 11, -12);
    elsif (x=73) then return to_sfixed(0.013698630137, 11, -12);
    elsif (x=74) then return to_sfixed(0.013513513514, 11, -12);
    elsif (x=75) then return to_sfixed(0.013333333333, 11, -12);
    elsif (x=76) then return to_sfixed(0.013157894737, 11, -12);
    elsif (x=77) then return to_sfixed(0.012987012987, 11, -12);
    elsif (x=78) then return to_sfixed(0.012820512821, 11, -12);
    elsif (x=79) then return to_sfixed(0.012658227848, 11, -12);
    elsif (x=80) then return to_sfixed(0.012500000000, 11, -12);
    elsif (x=81) then return to_sfixed(0.012345679012, 11, -12);
    elsif (x=82) then return to_sfixed(0.012195121951, 11, -12);
    elsif (x=83) then return to_sfixed(0.012048192771, 11, -12);
    elsif (x=84) then return to_sfixed(0.011904761905, 11, -12);
    elsif (x=85) then return to_sfixed(0.011764705882, 11, -12);
    elsif (x=86) then return to_sfixed(0.011627906977, 11, -12);
    elsif (x=87) then return to_sfixed(0.011494252874, 11, -12);
    elsif (x=88) then return to_sfixed(0.011363636364, 11, -12);
    elsif (x=89) then return to_sfixed(0.011235955056, 11, -12);
    elsif (x=90) then return to_sfixed(0.011111111111, 11, -12);
    elsif (x=91) then return to_sfixed(0.010989010989, 11, -12);
    elsif (x=92) then return to_sfixed(0.010869565217, 11, -12);
    elsif (x=93) then return to_sfixed(0.010752688172, 11, -12);
    elsif (x=94) then return to_sfixed(0.010638297872, 11, -12);
    elsif (x=95) then return to_sfixed(0.010526315789, 11, -12);
    elsif (x=96) then return to_sfixed(0.010416666667, 11, -12);
    elsif (x=97) then return to_sfixed(0.010309278351, 11, -12);
    elsif (x=98) then return to_sfixed(0.010204081633, 11, -12);
    elsif (x=99) then return to_sfixed(0.010101010101, 11, -12);
    elsif (x=100) then return to_sfixed(0.010000000000, 11, -12);
    elsif (x=101) then return to_sfixed(0.009900990099, 11, -12);
    elsif (x=102) then return to_sfixed(0.009803921569, 11, -12);
    elsif (x=103) then return to_sfixed(0.009708737864, 11, -12);
    elsif (x=104) then return to_sfixed(0.009615384615, 11, -12);
    elsif (x=105) then return to_sfixed(0.009523809524, 11, -12);
    elsif (x=106) then return to_sfixed(0.009433962264, 11, -12);
    elsif (x=107) then return to_sfixed(0.009345794393, 11, -12);
    elsif (x=108) then return to_sfixed(0.009259259259, 11, -12);
    elsif (x=109) then return to_sfixed(0.009174311927, 11, -12);
    elsif (x=110) then return to_sfixed(0.009090909091, 11, -12);
    elsif (x=111) then return to_sfixed(0.009009009009, 11, -12);
    elsif (x=112) then return to_sfixed(0.008928571429, 11, -12);
    elsif (x=113) then return to_sfixed(0.008849557522, 11, -12);
    elsif (x=114) then return to_sfixed(0.008771929825, 11, -12);
    elsif (x=115) then return to_sfixed(0.008695652174, 11, -12);
    elsif (x=116) then return to_sfixed(0.008620689655, 11, -12);
    elsif (x=117) then return to_sfixed(0.008547008547, 11, -12);
    elsif (x=118) then return to_sfixed(0.008474576271, 11, -12);
    elsif (x=119) then return to_sfixed(0.008403361345, 11, -12);
    elsif (x=120) then return to_sfixed(0.008333333333, 11, -12);
    elsif (x=121) then return to_sfixed(0.008264462810, 11, -12);
    elsif (x=122) then return to_sfixed(0.008196721311, 11, -12);
    elsif (x=123) then return to_sfixed(0.008130081301, 11, -12);
    elsif (x=124) then return to_sfixed(0.008064516129, 11, -12);
    elsif (x=125) then return to_sfixed(0.008000000000, 11, -12);
    elsif (x=126) then return to_sfixed(0.007936507937, 11, -12);
    elsif (x=127) then return to_sfixed(0.007874015748, 11, -12);
    elsif (x=128) then return to_sfixed(0.007812500000, 11, -12);
    elsif (x=129) then return to_sfixed(0.007751937984, 11, -12);
    elsif (x=130) then return to_sfixed(0.007692307692, 11, -12);
    elsif (x=131) then return to_sfixed(0.007633587786, 11, -12);
    elsif (x=132) then return to_sfixed(0.007575757576, 11, -12);
    elsif (x=133) then return to_sfixed(0.007518796992, 11, -12);
    elsif (x=134) then return to_sfixed(0.007462686567, 11, -12);
    elsif (x=135) then return to_sfixed(0.007407407407, 11, -12);
    elsif (x=136) then return to_sfixed(0.007352941176, 11, -12);
    elsif (x=137) then return to_sfixed(0.007299270073, 11, -12);
    elsif (x=138) then return to_sfixed(0.007246376812, 11, -12);
    elsif (x=139) then return to_sfixed(0.007194244604, 11, -12);
    elsif (x=140) then return to_sfixed(0.007142857143, 11, -12);
    elsif (x=141) then return to_sfixed(0.007092198582, 11, -12);
    elsif (x=142) then return to_sfixed(0.007042253521, 11, -12);
    elsif (x=143) then return to_sfixed(0.006993006993, 11, -12);
    elsif (x=144) then return to_sfixed(0.006944444444, 11, -12);
    elsif (x=145) then return to_sfixed(0.006896551724, 11, -12);
    elsif (x=146) then return to_sfixed(0.006849315068, 11, -12);
    elsif (x=147) then return to_sfixed(0.006802721088, 11, -12);
    elsif (x=148) then return to_sfixed(0.006756756757, 11, -12);
    elsif (x=149) then return to_sfixed(0.006711409396, 11, -12);
    elsif (x=150) then return to_sfixed(0.006666666667, 11, -12);
    elsif (x=151) then return to_sfixed(0.006622516556, 11, -12);
    elsif (x=152) then return to_sfixed(0.006578947368, 11, -12);
    elsif (x=153) then return to_sfixed(0.006535947712, 11, -12);
    elsif (x=154) then return to_sfixed(0.006493506494, 11, -12);
    elsif (x=155) then return to_sfixed(0.006451612903, 11, -12);
    elsif (x=156) then return to_sfixed(0.006410256410, 11, -12);
    elsif (x=157) then return to_sfixed(0.006369426752, 11, -12);
    elsif (x=158) then return to_sfixed(0.006329113924, 11, -12);
    elsif (x=159) then return to_sfixed(0.006289308176, 11, -12);
    elsif (x=160) then return to_sfixed(0.006250000000, 11, -12);
    elsif (x=161) then return to_sfixed(0.006211180124, 11, -12);
    elsif (x=162) then return to_sfixed(0.006172839506, 11, -12);
    elsif (x=163) then return to_sfixed(0.006134969325, 11, -12);
    elsif (x=164) then return to_sfixed(0.006097560976, 11, -12);
    elsif (x=165) then return to_sfixed(0.006060606061, 11, -12);
    elsif (x=166) then return to_sfixed(0.006024096386, 11, -12);
    elsif (x=167) then return to_sfixed(0.005988023952, 11, -12);
    elsif (x=168) then return to_sfixed(0.005952380952, 11, -12);
    elsif (x=169) then return to_sfixed(0.005917159763, 11, -12);
    elsif (x=170) then return to_sfixed(0.005882352941, 11, -12);
    elsif (x=171) then return to_sfixed(0.005847953216, 11, -12);
    elsif (x=172) then return to_sfixed(0.005813953488, 11, -12);
    elsif (x=173) then return to_sfixed(0.005780346821, 11, -12);
    elsif (x=174) then return to_sfixed(0.005747126437, 11, -12);
    elsif (x=175) then return to_sfixed(0.005714285714, 11, -12);
    elsif (x=176) then return to_sfixed(0.005681818182, 11, -12);
    elsif (x=177) then return to_sfixed(0.005649717514, 11, -12);
    elsif (x=178) then return to_sfixed(0.005617977528, 11, -12);
    elsif (x=179) then return to_sfixed(0.005586592179, 11, -12);
    elsif (x=180) then return to_sfixed(0.005555555556, 11, -12);
    elsif (x=181) then return to_sfixed(0.005524861878, 11, -12);
    elsif (x=182) then return to_sfixed(0.005494505495, 11, -12);
    elsif (x=183) then return to_sfixed(0.005464480874, 11, -12);
    elsif (x=184) then return to_sfixed(0.005434782609, 11, -12);
    elsif (x=185) then return to_sfixed(0.005405405405, 11, -12);
    elsif (x=186) then return to_sfixed(0.005376344086, 11, -12);
    elsif (x=187) then return to_sfixed(0.005347593583, 11, -12);
    elsif (x=188) then return to_sfixed(0.005319148936, 11, -12);
    elsif (x=189) then return to_sfixed(0.005291005291, 11, -12);
    elsif (x=190) then return to_sfixed(0.005263157895, 11, -12);
    elsif (x=191) then return to_sfixed(0.005235602094, 11, -12);
    elsif (x=192) then return to_sfixed(0.005208333333, 11, -12);
    elsif (x=193) then return to_sfixed(0.005181347150, 11, -12);
    elsif (x=194) then return to_sfixed(0.005154639175, 11, -12);
    elsif (x=195) then return to_sfixed(0.005128205128, 11, -12);
    elsif (x=196) then return to_sfixed(0.005102040816, 11, -12);
    elsif (x=197) then return to_sfixed(0.005076142132, 11, -12);
    elsif (x=198) then return to_sfixed(0.005050505051, 11, -12);
    elsif (x=199) then return to_sfixed(0.005025125628, 11, -12);
    elsif (x=200) then return to_sfixed(0.005000000000, 11, -12);
    elsif (x=201) then return to_sfixed(0.004975124378, 11, -12);
    elsif (x=202) then return to_sfixed(0.004950495050, 11, -12);
    elsif (x=203) then return to_sfixed(0.004926108374, 11, -12);
    elsif (x=204) then return to_sfixed(0.004901960784, 11, -12);
    elsif (x=205) then return to_sfixed(0.004878048780, 11, -12);
    elsif (x=206) then return to_sfixed(0.004854368932, 11, -12);
    elsif (x=207) then return to_sfixed(0.004830917874, 11, -12);
    elsif (x=208) then return to_sfixed(0.004807692308, 11, -12);
    elsif (x=209) then return to_sfixed(0.004784688995, 11, -12);
    elsif (x=210) then return to_sfixed(0.004761904762, 11, -12);
    elsif (x=211) then return to_sfixed(0.004739336493, 11, -12);
    elsif (x=212) then return to_sfixed(0.004716981132, 11, -12);
    elsif (x=213) then return to_sfixed(0.004694835681, 11, -12);
    elsif (x=214) then return to_sfixed(0.004672897196, 11, -12);
    elsif (x=215) then return to_sfixed(0.004651162791, 11, -12);
    elsif (x=216) then return to_sfixed(0.004629629630, 11, -12);
    elsif (x=217) then return to_sfixed(0.004608294931, 11, -12);
    elsif (x=218) then return to_sfixed(0.004587155963, 11, -12);
    elsif (x=219) then return to_sfixed(0.004566210046, 11, -12);
    elsif (x=220) then return to_sfixed(0.004545454545, 11, -12);
    elsif (x=221) then return to_sfixed(0.004524886878, 11, -12);
    elsif (x=222) then return to_sfixed(0.004504504505, 11, -12);
    elsif (x=223) then return to_sfixed(0.004484304933, 11, -12);
    elsif (x=224) then return to_sfixed(0.004464285714, 11, -12);
    elsif (x=225) then return to_sfixed(0.004444444444, 11, -12);
    elsif (x=226) then return to_sfixed(0.004424778761, 11, -12);
    elsif (x=227) then return to_sfixed(0.004405286344, 11, -12);
    elsif (x=228) then return to_sfixed(0.004385964912, 11, -12);
    elsif (x=229) then return to_sfixed(0.004366812227, 11, -12);
    elsif (x=230) then return to_sfixed(0.004347826087, 11, -12);
    elsif (x=231) then return to_sfixed(0.004329004329, 11, -12);
    elsif (x=232) then return to_sfixed(0.004310344828, 11, -12);
    elsif (x=233) then return to_sfixed(0.004291845494, 11, -12);
    elsif (x=234) then return to_sfixed(0.004273504274, 11, -12);
    elsif (x=235) then return to_sfixed(0.004255319149, 11, -12);
    elsif (x=236) then return to_sfixed(0.004237288136, 11, -12);
    elsif (x=237) then return to_sfixed(0.004219409283, 11, -12);
    elsif (x=238) then return to_sfixed(0.004201680672, 11, -12);
    elsif (x=239) then return to_sfixed(0.004184100418, 11, -12);
    elsif (x=240) then return to_sfixed(0.004166666667, 11, -12);
    elsif (x=241) then return to_sfixed(0.004149377593, 11, -12);
    elsif (x=242) then return to_sfixed(0.004132231405, 11, -12);
    elsif (x=243) then return to_sfixed(0.004115226337, 11, -12);
    elsif (x=244) then return to_sfixed(0.004098360656, 11, -12);
    elsif (x=245) then return to_sfixed(0.004081632653, 11, -12);
    elsif (x=246) then return to_sfixed(0.004065040650, 11, -12);
    elsif (x=247) then return to_sfixed(0.004048582996, 11, -12);
    elsif (x=248) then return to_sfixed(0.004032258065, 11, -12);
    elsif (x=249) then return to_sfixed(0.004016064257, 11, -12);
    elsif (x=250) then return to_sfixed(0.004000000000, 11, -12);
    elsif (x=251) then return to_sfixed(0.003984063745, 11, -12);
    elsif (x=252) then return to_sfixed(0.003968253968, 11, -12);
    elsif (x=253) then return to_sfixed(0.003952569170, 11, -12);
    elsif (x=254) then return to_sfixed(0.003937007874, 11, -12);
    elsif (x=255) then return to_sfixed(0.003921568627, 11, -12);
    elsif (x=256) then return to_sfixed(0.003906250000, 11, -12);
    elsif (x=257) then return to_sfixed(0.003891050584, 11, -12);
    elsif (x=258) then return to_sfixed(0.003875968992, 11, -12);
    elsif (x=259) then return to_sfixed(0.003861003861, 11, -12);
    elsif (x=260) then return to_sfixed(0.003846153846, 11, -12);
    elsif (x=261) then return to_sfixed(0.003831417625, 11, -12);
    elsif (x=262) then return to_sfixed(0.003816793893, 11, -12);
    elsif (x=263) then return to_sfixed(0.003802281369, 11, -12);
    elsif (x=264) then return to_sfixed(0.003787878788, 11, -12);
    elsif (x=265) then return to_sfixed(0.003773584906, 11, -12);
    elsif (x=266) then return to_sfixed(0.003759398496, 11, -12);
    elsif (x=267) then return to_sfixed(0.003745318352, 11, -12);
    elsif (x=268) then return to_sfixed(0.003731343284, 11, -12);
    elsif (x=269) then return to_sfixed(0.003717472119, 11, -12);
    elsif (x=270) then return to_sfixed(0.003703703704, 11, -12);
    elsif (x=271) then return to_sfixed(0.003690036900, 11, -12);
    elsif (x=272) then return to_sfixed(0.003676470588, 11, -12);
    elsif (x=273) then return to_sfixed(0.003663003663, 11, -12);
    elsif (x=274) then return to_sfixed(0.003649635036, 11, -12);
    elsif (x=275) then return to_sfixed(0.003636363636, 11, -12);
    elsif (x=276) then return to_sfixed(0.003623188406, 11, -12);
    elsif (x=277) then return to_sfixed(0.003610108303, 11, -12);
    elsif (x=278) then return to_sfixed(0.003597122302, 11, -12);
    elsif (x=279) then return to_sfixed(0.003584229391, 11, -12);
    elsif (x=280) then return to_sfixed(0.003571428571, 11, -12);
    elsif (x=281) then return to_sfixed(0.003558718861, 11, -12);
    elsif (x=282) then return to_sfixed(0.003546099291, 11, -12);
    elsif (x=283) then return to_sfixed(0.003533568905, 11, -12);
    elsif (x=284) then return to_sfixed(0.003521126761, 11, -12);
    elsif (x=285) then return to_sfixed(0.003508771930, 11, -12);
    elsif (x=286) then return to_sfixed(0.003496503497, 11, -12);
    elsif (x=287) then return to_sfixed(0.003484320557, 11, -12);
    elsif (x=288) then return to_sfixed(0.003472222222, 11, -12);
    elsif (x=289) then return to_sfixed(0.003460207612, 11, -12);
    elsif (x=290) then return to_sfixed(0.003448275862, 11, -12);
    elsif (x=291) then return to_sfixed(0.003436426117, 11, -12);
    elsif (x=292) then return to_sfixed(0.003424657534, 11, -12);
    elsif (x=293) then return to_sfixed(0.003412969283, 11, -12);
    elsif (x=294) then return to_sfixed(0.003401360544, 11, -12);
    elsif (x=295) then return to_sfixed(0.003389830508, 11, -12);
    elsif (x=296) then return to_sfixed(0.003378378378, 11, -12);
    elsif (x=297) then return to_sfixed(0.003367003367, 11, -12);
    elsif (x=298) then return to_sfixed(0.003355704698, 11, -12);
    elsif (x=299) then return to_sfixed(0.003344481605, 11, -12);
    elsif (x=300) then return to_sfixed(0.003333333333, 11, -12);
    elsif (x=301) then return to_sfixed(0.003322259136, 11, -12);
    elsif (x=302) then return to_sfixed(0.003311258278, 11, -12);
    elsif (x=303) then return to_sfixed(0.003300330033, 11, -12);
    elsif (x=304) then return to_sfixed(0.003289473684, 11, -12);
    elsif (x=305) then return to_sfixed(0.003278688525, 11, -12);
    elsif (x=306) then return to_sfixed(0.003267973856, 11, -12);
    elsif (x=307) then return to_sfixed(0.003257328990, 11, -12);
    elsif (x=308) then return to_sfixed(0.003246753247, 11, -12);
    elsif (x=309) then return to_sfixed(0.003236245955, 11, -12);
    elsif (x=310) then return to_sfixed(0.003225806452, 11, -12);
    elsif (x=311) then return to_sfixed(0.003215434084, 11, -12);
    elsif (x=312) then return to_sfixed(0.003205128205, 11, -12);
    elsif (x=313) then return to_sfixed(0.003194888179, 11, -12);
    elsif (x=314) then return to_sfixed(0.003184713376, 11, -12);
    elsif (x=315) then return to_sfixed(0.003174603175, 11, -12);
    elsif (x=316) then return to_sfixed(0.003164556962, 11, -12);
    elsif (x=317) then return to_sfixed(0.003154574132, 11, -12);
    elsif (x=318) then return to_sfixed(0.003144654088, 11, -12);
    elsif (x=319) then return to_sfixed(0.003134796238, 11, -12);
    elsif (x=320) then return to_sfixed(0.003125000000, 11, -12);
    elsif (x=321) then return to_sfixed(0.003115264798, 11, -12);
    elsif (x=322) then return to_sfixed(0.003105590062, 11, -12);
    elsif (x=323) then return to_sfixed(0.003095975232, 11, -12);
    elsif (x=324) then return to_sfixed(0.003086419753, 11, -12);
    elsif (x=325) then return to_sfixed(0.003076923077, 11, -12);
    elsif (x=326) then return to_sfixed(0.003067484663, 11, -12);
    elsif (x=327) then return to_sfixed(0.003058103976, 11, -12);
    elsif (x=328) then return to_sfixed(0.003048780488, 11, -12);
    elsif (x=329) then return to_sfixed(0.003039513678, 11, -12);
    elsif (x=330) then return to_sfixed(0.003030303030, 11, -12);
    elsif (x=331) then return to_sfixed(0.003021148036, 11, -12);
    elsif (x=332) then return to_sfixed(0.003012048193, 11, -12);
    elsif (x=333) then return to_sfixed(0.003003003003, 11, -12);
    elsif (x=334) then return to_sfixed(0.002994011976, 11, -12);
    elsif (x=335) then return to_sfixed(0.002985074627, 11, -12);
    elsif (x=336) then return to_sfixed(0.002976190476, 11, -12);
    elsif (x=337) then return to_sfixed(0.002967359050, 11, -12);
    elsif (x=338) then return to_sfixed(0.002958579882, 11, -12);
    elsif (x=339) then return to_sfixed(0.002949852507, 11, -12);
    elsif (x=340) then return to_sfixed(0.002941176471, 11, -12);
    elsif (x=341) then return to_sfixed(0.002932551320, 11, -12);
    elsif (x=342) then return to_sfixed(0.002923976608, 11, -12);
    elsif (x=343) then return to_sfixed(0.002915451895, 11, -12);
    elsif (x=344) then return to_sfixed(0.002906976744, 11, -12);
    elsif (x=345) then return to_sfixed(0.002898550725, 11, -12);
    elsif (x=346) then return to_sfixed(0.002890173410, 11, -12);
    elsif (x=347) then return to_sfixed(0.002881844380, 11, -12);
    elsif (x=348) then return to_sfixed(0.002873563218, 11, -12);
    elsif (x=349) then return to_sfixed(0.002865329513, 11, -12);
    elsif (x=350) then return to_sfixed(0.002857142857, 11, -12);
    elsif (x=351) then return to_sfixed(0.002849002849, 11, -12);
    elsif (x=352) then return to_sfixed(0.002840909091, 11, -12);
    elsif (x=353) then return to_sfixed(0.002832861190, 11, -12);
    elsif (x=354) then return to_sfixed(0.002824858757, 11, -12);
    elsif (x=355) then return to_sfixed(0.002816901408, 11, -12);
    elsif (x=356) then return to_sfixed(0.002808988764, 11, -12);
    elsif (x=357) then return to_sfixed(0.002801120448, 11, -12);
    elsif (x=358) then return to_sfixed(0.002793296089, 11, -12);
    elsif (x=359) then return to_sfixed(0.002785515320, 11, -12);
    elsif (x=360) then return to_sfixed(0.002777777778, 11, -12);
    elsif (x=361) then return to_sfixed(0.002770083102, 11, -12);
    elsif (x=362) then return to_sfixed(0.002762430939, 11, -12);
    elsif (x=363) then return to_sfixed(0.002754820937, 11, -12);
    elsif (x=364) then return to_sfixed(0.002747252747, 11, -12);
    elsif (x=365) then return to_sfixed(0.002739726027, 11, -12);
    elsif (x=366) then return to_sfixed(0.002732240437, 11, -12);
    elsif (x=367) then return to_sfixed(0.002724795640, 11, -12);
    elsif (x=368) then return to_sfixed(0.002717391304, 11, -12);
    elsif (x=369) then return to_sfixed(0.002710027100, 11, -12);
    elsif (x=370) then return to_sfixed(0.002702702703, 11, -12);
    elsif (x=371) then return to_sfixed(0.002695417790, 11, -12);
    elsif (x=372) then return to_sfixed(0.002688172043, 11, -12);
    elsif (x=373) then return to_sfixed(0.002680965147, 11, -12);
    elsif (x=374) then return to_sfixed(0.002673796791, 11, -12);
    elsif (x=375) then return to_sfixed(0.002666666667, 11, -12);
    elsif (x=376) then return to_sfixed(0.002659574468, 11, -12);
    elsif (x=377) then return to_sfixed(0.002652519894, 11, -12);
    elsif (x=378) then return to_sfixed(0.002645502646, 11, -12);
    elsif (x=379) then return to_sfixed(0.002638522427, 11, -12);
    elsif (x=380) then return to_sfixed(0.002631578947, 11, -12);
    elsif (x=381) then return to_sfixed(0.002624671916, 11, -12);
    elsif (x=382) then return to_sfixed(0.002617801047, 11, -12);
    elsif (x=383) then return to_sfixed(0.002610966057, 11, -12);
    elsif (x=384) then return to_sfixed(0.002604166667, 11, -12);
    elsif (x=385) then return to_sfixed(0.002597402597, 11, -12);
    elsif (x=386) then return to_sfixed(0.002590673575, 11, -12);
    elsif (x=387) then return to_sfixed(0.002583979328, 11, -12);
    elsif (x=388) then return to_sfixed(0.002577319588, 11, -12);
    elsif (x=389) then return to_sfixed(0.002570694087, 11, -12);
    elsif (x=390) then return to_sfixed(0.002564102564, 11, -12);
    elsif (x=391) then return to_sfixed(0.002557544757, 11, -12);
    elsif (x=392) then return to_sfixed(0.002551020408, 11, -12);
    elsif (x=393) then return to_sfixed(0.002544529262, 11, -12);
    elsif (x=394) then return to_sfixed(0.002538071066, 11, -12);
    elsif (x=395) then return to_sfixed(0.002531645570, 11, -12);
    elsif (x=396) then return to_sfixed(0.002525252525, 11, -12);
    elsif (x=397) then return to_sfixed(0.002518891688, 11, -12);
    elsif (x=398) then return to_sfixed(0.002512562814, 11, -12);
    elsif (x=399) then return to_sfixed(0.002506265664, 11, -12);
    elsif (x=400) then return to_sfixed(0.002500000000, 11, -12);
    elsif (x=401) then return to_sfixed(0.002493765586, 11, -12);
    elsif (x=402) then return to_sfixed(0.002487562189, 11, -12);
    elsif (x=403) then return to_sfixed(0.002481389578, 11, -12);
    elsif (x=404) then return to_sfixed(0.002475247525, 11, -12);
    elsif (x=405) then return to_sfixed(0.002469135802, 11, -12);
    elsif (x=406) then return to_sfixed(0.002463054187, 11, -12);
    elsif (x=407) then return to_sfixed(0.002457002457, 11, -12);
    elsif (x=408) then return to_sfixed(0.002450980392, 11, -12);
    elsif (x=409) then return to_sfixed(0.002444987775, 11, -12);
    elsif (x=410) then return to_sfixed(0.002439024390, 11, -12);
    elsif (x=411) then return to_sfixed(0.002433090024, 11, -12);
    elsif (x=412) then return to_sfixed(0.002427184466, 11, -12);
    elsif (x=413) then return to_sfixed(0.002421307506, 11, -12);
    elsif (x=414) then return to_sfixed(0.002415458937, 11, -12);
    elsif (x=415) then return to_sfixed(0.002409638554, 11, -12);
    elsif (x=416) then return to_sfixed(0.002403846154, 11, -12);
    elsif (x=417) then return to_sfixed(0.002398081535, 11, -12);
    elsif (x=418) then return to_sfixed(0.002392344498, 11, -12);
    elsif (x=419) then return to_sfixed(0.002386634845, 11, -12);
    elsif (x=420) then return to_sfixed(0.002380952381, 11, -12);
    elsif (x=421) then return to_sfixed(0.002375296912, 11, -12);
    elsif (x=422) then return to_sfixed(0.002369668246, 11, -12);
    elsif (x=423) then return to_sfixed(0.002364066194, 11, -12);
    elsif (x=424) then return to_sfixed(0.002358490566, 11, -12);
    elsif (x=425) then return to_sfixed(0.002352941176, 11, -12);
    elsif (x=426) then return to_sfixed(0.002347417840, 11, -12);
    elsif (x=427) then return to_sfixed(0.002341920375, 11, -12);
    elsif (x=428) then return to_sfixed(0.002336448598, 11, -12);
    elsif (x=429) then return to_sfixed(0.002331002331, 11, -12);
    elsif (x=430) then return to_sfixed(0.002325581395, 11, -12);
    elsif (x=431) then return to_sfixed(0.002320185615, 11, -12);
    elsif (x=432) then return to_sfixed(0.002314814815, 11, -12);
    elsif (x=433) then return to_sfixed(0.002309468822, 11, -12);
    elsif (x=434) then return to_sfixed(0.002304147465, 11, -12);
    elsif (x=435) then return to_sfixed(0.002298850575, 11, -12);
    elsif (x=436) then return to_sfixed(0.002293577982, 11, -12);
    elsif (x=437) then return to_sfixed(0.002288329519, 11, -12);
    elsif (x=438) then return to_sfixed(0.002283105023, 11, -12);
    elsif (x=439) then return to_sfixed(0.002277904328, 11, -12);
    elsif (x=440) then return to_sfixed(0.002272727273, 11, -12);
    elsif (x=441) then return to_sfixed(0.002267573696, 11, -12);
    elsif (x=442) then return to_sfixed(0.002262443439, 11, -12);
    elsif (x=443) then return to_sfixed(0.002257336343, 11, -12);
    elsif (x=444) then return to_sfixed(0.002252252252, 11, -12);
    elsif (x=445) then return to_sfixed(0.002247191011, 11, -12);
    elsif (x=446) then return to_sfixed(0.002242152466, 11, -12);
    elsif (x=447) then return to_sfixed(0.002237136465, 11, -12);
    elsif (x=448) then return to_sfixed(0.002232142857, 11, -12);
    elsif (x=449) then return to_sfixed(0.002227171492, 11, -12);
    elsif (x=450) then return to_sfixed(0.002222222222, 11, -12);
    elsif (x=451) then return to_sfixed(0.002217294900, 11, -12);
    elsif (x=452) then return to_sfixed(0.002212389381, 11, -12);
    elsif (x=453) then return to_sfixed(0.002207505519, 11, -12);
    elsif (x=454) then return to_sfixed(0.002202643172, 11, -12);
    elsif (x=455) then return to_sfixed(0.002197802198, 11, -12);
    elsif (x=456) then return to_sfixed(0.002192982456, 11, -12);
    elsif (x=457) then return to_sfixed(0.002188183807, 11, -12);
    elsif (x=458) then return to_sfixed(0.002183406114, 11, -12);
    elsif (x=459) then return to_sfixed(0.002178649237, 11, -12);
    elsif (x=460) then return to_sfixed(0.002173913043, 11, -12);
    elsif (x=461) then return to_sfixed(0.002169197397, 11, -12);
    elsif (x=462) then return to_sfixed(0.002164502165, 11, -12);
    elsif (x=463) then return to_sfixed(0.002159827214, 11, -12);
    elsif (x=464) then return to_sfixed(0.002155172414, 11, -12);
    elsif (x=465) then return to_sfixed(0.002150537634, 11, -12);
    elsif (x=466) then return to_sfixed(0.002145922747, 11, -12);
    elsif (x=467) then return to_sfixed(0.002141327623, 11, -12);
    elsif (x=468) then return to_sfixed(0.002136752137, 11, -12);
    elsif (x=469) then return to_sfixed(0.002132196162, 11, -12);
    elsif (x=470) then return to_sfixed(0.002127659574, 11, -12);
    elsif (x=471) then return to_sfixed(0.002123142251, 11, -12);
    elsif (x=472) then return to_sfixed(0.002118644068, 11, -12);
    elsif (x=473) then return to_sfixed(0.002114164905, 11, -12);
    elsif (x=474) then return to_sfixed(0.002109704641, 11, -12);
    elsif (x=475) then return to_sfixed(0.002105263158, 11, -12);
    elsif (x=476) then return to_sfixed(0.002100840336, 11, -12);
    elsif (x=477) then return to_sfixed(0.002096436059, 11, -12);
    elsif (x=478) then return to_sfixed(0.002092050209, 11, -12);
    elsif (x=479) then return to_sfixed(0.002087682672, 11, -12);
    elsif (x=480) then return to_sfixed(0.002083333333, 11, -12);
    elsif (x=481) then return to_sfixed(0.002079002079, 11, -12);
    elsif (x=482) then return to_sfixed(0.002074688797, 11, -12);
    elsif (x=483) then return to_sfixed(0.002070393375, 11, -12);
    elsif (x=484) then return to_sfixed(0.002066115702, 11, -12);
    elsif (x=485) then return to_sfixed(0.002061855670, 11, -12);
    elsif (x=486) then return to_sfixed(0.002057613169, 11, -12);
    elsif (x=487) then return to_sfixed(0.002053388090, 11, -12);
    elsif (x=488) then return to_sfixed(0.002049180328, 11, -12);
    elsif (x=489) then return to_sfixed(0.002044989775, 11, -12);
    elsif (x=490) then return to_sfixed(0.002040816327, 11, -12);
    elsif (x=491) then return to_sfixed(0.002036659878, 11, -12);
    elsif (x=492) then return to_sfixed(0.002032520325, 11, -12);
    elsif (x=493) then return to_sfixed(0.002028397566, 11, -12);
    elsif (x=494) then return to_sfixed(0.002024291498, 11, -12);
    elsif (x=495) then return to_sfixed(0.002020202020, 11, -12);
    elsif (x=496) then return to_sfixed(0.002016129032, 11, -12);
    elsif (x=497) then return to_sfixed(0.002012072435, 11, -12);
    elsif (x=498) then return to_sfixed(0.002008032129, 11, -12);
    elsif (x=499) then return to_sfixed(0.002004008016, 11, -12);
    elsif (x=500) then return to_sfixed(0.002000000000, 11, -12);
    elsif (x=501) then return to_sfixed(0.001996007984, 11, -12);
    elsif (x=502) then return to_sfixed(0.001992031873, 11, -12);
    elsif (x=503) then return to_sfixed(0.001988071571, 11, -12);
    elsif (x=504) then return to_sfixed(0.001984126984, 11, -12);
    elsif (x=505) then return to_sfixed(0.001980198020, 11, -12);
    elsif (x=506) then return to_sfixed(0.001976284585, 11, -12);
    elsif (x=507) then return to_sfixed(0.001972386588, 11, -12);
    elsif (x=508) then return to_sfixed(0.001968503937, 11, -12);
    elsif (x=509) then return to_sfixed(0.001964636542, 11, -12);
    elsif (x=510) then return to_sfixed(0.001960784314, 11, -12);
    elsif (x=511) then return to_sfixed(0.001956947162, 11, -12);
    elsif (x=512) then return to_sfixed(0.001953125000, 11, -12);
    elsif (x=513) then return to_sfixed(0.001949317739, 11, -12);
    elsif (x=514) then return to_sfixed(0.001945525292, 11, -12);
    elsif (x=515) then return to_sfixed(0.001941747573, 11, -12);
    elsif (x=516) then return to_sfixed(0.001937984496, 11, -12);
    elsif (x=517) then return to_sfixed(0.001934235977, 11, -12);
    elsif (x=518) then return to_sfixed(0.001930501931, 11, -12);
    elsif (x=519) then return to_sfixed(0.001926782274, 11, -12);
    elsif (x=520) then return to_sfixed(0.001923076923, 11, -12);
    elsif (x=521) then return to_sfixed(0.001919385797, 11, -12);
    elsif (x=522) then return to_sfixed(0.001915708812, 11, -12);
    elsif (x=523) then return to_sfixed(0.001912045889, 11, -12);
    elsif (x=524) then return to_sfixed(0.001908396947, 11, -12);
    elsif (x=525) then return to_sfixed(0.001904761905, 11, -12);
    elsif (x=526) then return to_sfixed(0.001901140684, 11, -12);
    elsif (x=527) then return to_sfixed(0.001897533207, 11, -12);
    elsif (x=528) then return to_sfixed(0.001893939394, 11, -12);
    elsif (x=529) then return to_sfixed(0.001890359168, 11, -12);
    elsif (x=530) then return to_sfixed(0.001886792453, 11, -12);
    elsif (x=531) then return to_sfixed(0.001883239171, 11, -12);
    elsif (x=532) then return to_sfixed(0.001879699248, 11, -12);
    elsif (x=533) then return to_sfixed(0.001876172608, 11, -12);
    elsif (x=534) then return to_sfixed(0.001872659176, 11, -12);
    elsif (x=535) then return to_sfixed(0.001869158879, 11, -12);
    elsif (x=536) then return to_sfixed(0.001865671642, 11, -12);
    elsif (x=537) then return to_sfixed(0.001862197393, 11, -12);
    elsif (x=538) then return to_sfixed(0.001858736059, 11, -12);
    elsif (x=539) then return to_sfixed(0.001855287570, 11, -12);
    elsif (x=540) then return to_sfixed(0.001851851852, 11, -12);
    elsif (x=541) then return to_sfixed(0.001848428835, 11, -12);
    elsif (x=542) then return to_sfixed(0.001845018450, 11, -12);
    elsif (x=543) then return to_sfixed(0.001841620626, 11, -12);
    elsif (x=544) then return to_sfixed(0.001838235294, 11, -12);
    elsif (x=545) then return to_sfixed(0.001834862385, 11, -12);
    elsif (x=546) then return to_sfixed(0.001831501832, 11, -12);
    elsif (x=547) then return to_sfixed(0.001828153565, 11, -12);
    elsif (x=548) then return to_sfixed(0.001824817518, 11, -12);
    elsif (x=549) then return to_sfixed(0.001821493625, 11, -12);
    elsif (x=550) then return to_sfixed(0.001818181818, 11, -12);
    elsif (x=551) then return to_sfixed(0.001814882033, 11, -12);
    elsif (x=552) then return to_sfixed(0.001811594203, 11, -12);
    elsif (x=553) then return to_sfixed(0.001808318264, 11, -12);
    elsif (x=554) then return to_sfixed(0.001805054152, 11, -12);
    elsif (x=555) then return to_sfixed(0.001801801802, 11, -12);
    elsif (x=556) then return to_sfixed(0.001798561151, 11, -12);
    elsif (x=557) then return to_sfixed(0.001795332136, 11, -12);
    elsif (x=558) then return to_sfixed(0.001792114695, 11, -12);
    elsif (x=559) then return to_sfixed(0.001788908766, 11, -12);
    elsif (x=560) then return to_sfixed(0.001785714286, 11, -12);
    elsif (x=561) then return to_sfixed(0.001782531194, 11, -12);
    elsif (x=562) then return to_sfixed(0.001779359431, 11, -12);
    elsif (x=563) then return to_sfixed(0.001776198934, 11, -12);
    elsif (x=564) then return to_sfixed(0.001773049645, 11, -12);
    elsif (x=565) then return to_sfixed(0.001769911504, 11, -12);
    elsif (x=566) then return to_sfixed(0.001766784452, 11, -12);
    elsif (x=567) then return to_sfixed(0.001763668430, 11, -12);
    elsif (x=568) then return to_sfixed(0.001760563380, 11, -12);
    elsif (x=569) then return to_sfixed(0.001757469244, 11, -12);
    elsif (x=570) then return to_sfixed(0.001754385965, 11, -12);
    elsif (x=571) then return to_sfixed(0.001751313485, 11, -12);
    elsif (x=572) then return to_sfixed(0.001748251748, 11, -12);
    elsif (x=573) then return to_sfixed(0.001745200698, 11, -12);
    elsif (x=574) then return to_sfixed(0.001742160279, 11, -12);
    elsif (x=575) then return to_sfixed(0.001739130435, 11, -12);
    elsif (x=576) then return to_sfixed(0.001736111111, 11, -12);
    elsif (x=577) then return to_sfixed(0.001733102253, 11, -12);
    elsif (x=578) then return to_sfixed(0.001730103806, 11, -12);
    elsif (x=579) then return to_sfixed(0.001727115717, 11, -12);
    elsif (x=580) then return to_sfixed(0.001724137931, 11, -12);
    elsif (x=581) then return to_sfixed(0.001721170396, 11, -12);
    elsif (x=582) then return to_sfixed(0.001718213058, 11, -12);
    elsif (x=583) then return to_sfixed(0.001715265866, 11, -12);
    elsif (x=584) then return to_sfixed(0.001712328767, 11, -12);
    elsif (x=585) then return to_sfixed(0.001709401709, 11, -12);
    elsif (x=586) then return to_sfixed(0.001706484642, 11, -12);
    elsif (x=587) then return to_sfixed(0.001703577513, 11, -12);
    elsif (x=588) then return to_sfixed(0.001700680272, 11, -12);
    elsif (x=589) then return to_sfixed(0.001697792869, 11, -12);
    elsif (x=590) then return to_sfixed(0.001694915254, 11, -12);
    elsif (x=591) then return to_sfixed(0.001692047377, 11, -12);
    elsif (x=592) then return to_sfixed(0.001689189189, 11, -12);
    elsif (x=593) then return to_sfixed(0.001686340641, 11, -12);
    elsif (x=594) then return to_sfixed(0.001683501684, 11, -12);
    elsif (x=595) then return to_sfixed(0.001680672269, 11, -12);
    elsif (x=596) then return to_sfixed(0.001677852349, 11, -12);
    elsif (x=597) then return to_sfixed(0.001675041876, 11, -12);
    elsif (x=598) then return to_sfixed(0.001672240803, 11, -12);
    elsif (x=599) then return to_sfixed(0.001669449082, 11, -12);
    elsif (x=600) then return to_sfixed(0.001666666667, 11, -12);
    elsif (x=601) then return to_sfixed(0.001663893511, 11, -12);
    elsif (x=602) then return to_sfixed(0.001661129568, 11, -12);
    elsif (x=603) then return to_sfixed(0.001658374793, 11, -12);
    elsif (x=604) then return to_sfixed(0.001655629139, 11, -12);
    elsif (x=605) then return to_sfixed(0.001652892562, 11, -12);
    elsif (x=606) then return to_sfixed(0.001650165017, 11, -12);
    elsif (x=607) then return to_sfixed(0.001647446458, 11, -12);
    elsif (x=608) then return to_sfixed(0.001644736842, 11, -12);
    elsif (x=609) then return to_sfixed(0.001642036125, 11, -12);
    elsif (x=610) then return to_sfixed(0.001639344262, 11, -12);
    elsif (x=611) then return to_sfixed(0.001636661211, 11, -12);
    elsif (x=612) then return to_sfixed(0.001633986928, 11, -12);
    elsif (x=613) then return to_sfixed(0.001631321370, 11, -12);
    elsif (x=614) then return to_sfixed(0.001628664495, 11, -12);
    elsif (x=615) then return to_sfixed(0.001626016260, 11, -12);
    elsif (x=616) then return to_sfixed(0.001623376623, 11, -12);
    elsif (x=617) then return to_sfixed(0.001620745543, 11, -12);
    elsif (x=618) then return to_sfixed(0.001618122977, 11, -12);
    elsif (x=619) then return to_sfixed(0.001615508885, 11, -12);
    elsif (x=620) then return to_sfixed(0.001612903226, 11, -12);
    elsif (x=621) then return to_sfixed(0.001610305958, 11, -12);
    elsif (x=622) then return to_sfixed(0.001607717042, 11, -12);
    elsif (x=623) then return to_sfixed(0.001605136437, 11, -12);
    elsif (x=624) then return to_sfixed(0.001602564103, 11, -12);
    elsif (x=625) then return to_sfixed(0.001600000000, 11, -12);
    elsif (x=626) then return to_sfixed(0.001597444089, 11, -12);
    elsif (x=627) then return to_sfixed(0.001594896332, 11, -12);
    elsif (x=628) then return to_sfixed(0.001592356688, 11, -12);
    elsif (x=629) then return to_sfixed(0.001589825119, 11, -12);
    elsif (x=630) then return to_sfixed(0.001587301587, 11, -12);
    end if;
  end;

end package body reciprocal_pkg;
