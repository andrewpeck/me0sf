
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

package sf_pkg is

  type partition_t is array (integer range 0 to 5) of std_logic_vector;

end package sf_pkg;
