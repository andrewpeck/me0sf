----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- ME0 Segment Finder Firmware
-- A. Peck, C. Grubb, J. Chismar
----------------------------------------------------------------------------------
-- Description:
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;



entity centroid_finder is

  generic(LENGTH : integer; NBITS : integer);

  port(

    clk : in std_logic;

    din : in std_logic_vector(LENGTH-1 downto 0);

    dout : out unsigned(NBITS-1 downto 0)

    );

end centroid_finder;



architecture behavioral of centroid_finder is

    signal index : natural range 0 to LENGTH;



begin

  gen_1 : if (length = 1) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din(0) is
         when '0' => index <= 0;
         when '1' => index <= 1;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_2 : if (length = 2) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "00" => index <= 0;
         when "01" => index <= 1;
         when "10" => index <= 2;
         when "11" => index <= 2;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_3 : if (length = 3) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "000" => index <= 0;
         when "001" => index <= 1;
         when "010" => index <= 2;
         when "011" => index <= 2;
         when "100" => index <= 3;
         when "101" => index <= 2;
         when "110" => index <= 2;
         when "111" => index <= 2;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_4 : if (length = 4) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "0000" => index <= 0;
         when "0001" => index <= 1;
         when "0010" => index <= 2;
         when "0011" => index <= 2;
         when "0100" => index <= 3;
         when "0101" => index <= 2;
         when "0110" => index <= 2;
         when "0111" => index <= 2;
         when "1000" => index <= 4;
         when "1001" => index <= 2;
         when "1010" => index <= 3;
         when "1011" => index <= 2;
         when "1100" => index <= 4;
         when "1101" => index <= 3;
         when "1110" => index <= 3;
         when "1111" => index <= 2;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_5 : if (length = 5) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "00000" => index <= 0;
         when "00001" => index <= 1;
         when "00010" => index <= 2;
         when "00011" => index <= 2;
         when "00100" => index <= 3;
         when "00101" => index <= 2;
         when "00110" => index <= 2;
         when "00111" => index <= 2;
         when "01000" => index <= 4;
         when "01001" => index <= 2;
         when "01010" => index <= 3;
         when "01011" => index <= 2;
         when "01100" => index <= 4;
         when "01101" => index <= 3;
         when "01110" => index <= 3;
         when "01111" => index <= 2;
         when "10000" => index <= 5;
         when "10001" => index <= 3;
         when "10010" => index <= 4;
         when "10011" => index <= 3;
         when "10100" => index <= 4;
         when "10101" => index <= 3;
         when "10110" => index <= 3;
         when "10111" => index <= 3;
         when "11000" => index <= 4;
         when "11001" => index <= 3;
         when "11010" => index <= 4;
         when "11011" => index <= 3;
         when "11100" => index <= 4;
         when "11101" => index <= 3;
         when "11110" => index <= 4;
         when "11111" => index <= 3;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_6 : if (length = 6) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "000000" => index <= 0;
         when "000001" => index <= 1;
         when "000010" => index <= 2;
         when "000011" => index <= 2;
         when "000100" => index <= 3;
         when "000101" => index <= 2;
         when "000110" => index <= 2;
         when "000111" => index <= 2;
         when "001000" => index <= 4;
         when "001001" => index <= 2;
         when "001010" => index <= 3;
         when "001011" => index <= 2;
         when "001100" => index <= 4;
         when "001101" => index <= 3;
         when "001110" => index <= 3;
         when "001111" => index <= 2;
         when "010000" => index <= 5;
         when "010001" => index <= 3;
         when "010010" => index <= 4;
         when "010011" => index <= 3;
         when "010100" => index <= 4;
         when "010101" => index <= 3;
         when "010110" => index <= 3;
         when "010111" => index <= 3;
         when "011000" => index <= 4;
         when "011001" => index <= 3;
         when "011010" => index <= 4;
         when "011011" => index <= 3;
         when "011100" => index <= 4;
         when "011101" => index <= 3;
         when "011110" => index <= 4;
         when "011111" => index <= 3;
         when "100000" => index <= 6;
         when "100001" => index <= 4;
         when "100010" => index <= 4;
         when "100011" => index <= 3;
         when "100100" => index <= 4;
         when "100101" => index <= 3;
         when "100110" => index <= 4;
         when "100111" => index <= 3;
         when "101000" => index <= 5;
         when "101001" => index <= 4;
         when "101010" => index <= 4;
         when "101011" => index <= 3;
         when "101100" => index <= 4;
         when "101101" => index <= 4;
         when "101110" => index <= 4;
         when "101111" => index <= 3;
         when "110000" => index <= 6;
         when "110001" => index <= 4;
         when "110010" => index <= 4;
         when "110011" => index <= 4;
         when "110100" => index <= 5;
         when "110101" => index <= 4;
         when "110110" => index <= 4;
         when "110111" => index <= 3;
         when "111000" => index <= 5;
         when "111001" => index <= 4;
         when "111010" => index <= 4;
         when "111011" => index <= 4;
         when "111100" => index <= 4;
         when "111101" => index <= 4;
         when "111110" => index <= 4;
         when "111111" => index <= 4;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_7 : if (length = 7) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "0000000" => index <= 0;
         when "0000001" => index <= 1;
         when "0000010" => index <= 2;
         when "0000011" => index <= 2;
         when "0000100" => index <= 3;
         when "0000101" => index <= 2;
         when "0000110" => index <= 2;
         when "0000111" => index <= 2;
         when "0001000" => index <= 4;
         when "0001001" => index <= 2;
         when "0001010" => index <= 3;
         when "0001011" => index <= 2;
         when "0001100" => index <= 4;
         when "0001101" => index <= 3;
         when "0001110" => index <= 3;
         when "0001111" => index <= 2;
         when "0010000" => index <= 5;
         when "0010001" => index <= 3;
         when "0010010" => index <= 4;
         when "0010011" => index <= 3;
         when "0010100" => index <= 4;
         when "0010101" => index <= 3;
         when "0010110" => index <= 3;
         when "0010111" => index <= 3;
         when "0011000" => index <= 4;
         when "0011001" => index <= 3;
         when "0011010" => index <= 4;
         when "0011011" => index <= 3;
         when "0011100" => index <= 4;
         when "0011101" => index <= 3;
         when "0011110" => index <= 4;
         when "0011111" => index <= 3;
         when "0100000" => index <= 6;
         when "0100001" => index <= 4;
         when "0100010" => index <= 4;
         when "0100011" => index <= 3;
         when "0100100" => index <= 4;
         when "0100101" => index <= 3;
         when "0100110" => index <= 4;
         when "0100111" => index <= 3;
         when "0101000" => index <= 5;
         when "0101001" => index <= 4;
         when "0101010" => index <= 4;
         when "0101011" => index <= 3;
         when "0101100" => index <= 4;
         when "0101101" => index <= 4;
         when "0101110" => index <= 4;
         when "0101111" => index <= 3;
         when "0110000" => index <= 6;
         when "0110001" => index <= 4;
         when "0110010" => index <= 4;
         when "0110011" => index <= 4;
         when "0110100" => index <= 5;
         when "0110101" => index <= 4;
         when "0110110" => index <= 4;
         when "0110111" => index <= 3;
         when "0111000" => index <= 5;
         when "0111001" => index <= 4;
         when "0111010" => index <= 4;
         when "0111011" => index <= 4;
         when "0111100" => index <= 4;
         when "0111101" => index <= 4;
         when "0111110" => index <= 4;
         when "0111111" => index <= 4;
         when "1000000" => index <= 7;
         when "1000001" => index <= 4;
         when "1000010" => index <= 4;
         when "1000011" => index <= 3;
         when "1000100" => index <= 5;
         when "1000101" => index <= 4;
         when "1000110" => index <= 4;
         when "1000111" => index <= 3;
         when "1001000" => index <= 6;
         when "1001001" => index <= 4;
         when "1001010" => index <= 4;
         when "1001011" => index <= 4;
         when "1001100" => index <= 5;
         when "1001101" => index <= 4;
         when "1001110" => index <= 4;
         when "1001111" => index <= 3;
         when "1010000" => index <= 6;
         when "1010001" => index <= 4;
         when "1010010" => index <= 5;
         when "1010011" => index <= 4;
         when "1010100" => index <= 5;
         when "1010101" => index <= 4;
         when "1010110" => index <= 4;
         when "1010111" => index <= 4;
         when "1011000" => index <= 5;
         when "1011001" => index <= 4;
         when "1011010" => index <= 4;
         when "1011011" => index <= 4;
         when "1011100" => index <= 5;
         when "1011101" => index <= 4;
         when "1011110" => index <= 4;
         when "1011111" => index <= 4;
         when "1100000" => index <= 6;
         when "1100001" => index <= 5;
         when "1100010" => index <= 5;
         when "1100011" => index <= 4;
         when "1100100" => index <= 5;
         when "1100101" => index <= 4;
         when "1100110" => index <= 4;
         when "1100111" => index <= 4;
         when "1101000" => index <= 6;
         when "1101001" => index <= 4;
         when "1101010" => index <= 5;
         when "1101011" => index <= 4;
         when "1101100" => index <= 5;
         when "1101101" => index <= 4;
         when "1101110" => index <= 4;
         when "1101111" => index <= 4;
         when "1110000" => index <= 6;
         when "1110001" => index <= 5;
         when "1110010" => index <= 5;
         when "1110011" => index <= 4;
         when "1110100" => index <= 5;
         when "1110101" => index <= 4;
         when "1110110" => index <= 5;
         when "1110111" => index <= 4;
         when "1111000" => index <= 6;
         when "1111001" => index <= 5;
         when "1111010" => index <= 5;
         when "1111011" => index <= 4;
         when "1111100" => index <= 5;
         when "1111101" => index <= 4;
         when "1111110" => index <= 4;
         when "1111111" => index <= 4;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_8 : if (length = 8) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "00000000" => index <= 0;
         when "00000001" => index <= 1;
         when "00000010" => index <= 2;
         when "00000011" => index <= 2;
         when "00000100" => index <= 3;
         when "00000101" => index <= 2;
         when "00000110" => index <= 2;
         when "00000111" => index <= 2;
         when "00001000" => index <= 4;
         when "00001001" => index <= 2;
         when "00001010" => index <= 3;
         when "00001011" => index <= 2;
         when "00001100" => index <= 4;
         when "00001101" => index <= 3;
         when "00001110" => index <= 3;
         when "00001111" => index <= 2;
         when "00010000" => index <= 5;
         when "00010001" => index <= 3;
         when "00010010" => index <= 4;
         when "00010011" => index <= 3;
         when "00010100" => index <= 4;
         when "00010101" => index <= 3;
         when "00010110" => index <= 3;
         when "00010111" => index <= 3;
         when "00011000" => index <= 4;
         when "00011001" => index <= 3;
         when "00011010" => index <= 4;
         when "00011011" => index <= 3;
         when "00011100" => index <= 4;
         when "00011101" => index <= 3;
         when "00011110" => index <= 4;
         when "00011111" => index <= 3;
         when "00100000" => index <= 6;
         when "00100001" => index <= 4;
         when "00100010" => index <= 4;
         when "00100011" => index <= 3;
         when "00100100" => index <= 4;
         when "00100101" => index <= 3;
         when "00100110" => index <= 4;
         when "00100111" => index <= 3;
         when "00101000" => index <= 5;
         when "00101001" => index <= 4;
         when "00101010" => index <= 4;
         when "00101011" => index <= 3;
         when "00101100" => index <= 4;
         when "00101101" => index <= 4;
         when "00101110" => index <= 4;
         when "00101111" => index <= 3;
         when "00110000" => index <= 6;
         when "00110001" => index <= 4;
         when "00110010" => index <= 4;
         when "00110011" => index <= 4;
         when "00110100" => index <= 5;
         when "00110101" => index <= 4;
         when "00110110" => index <= 4;
         when "00110111" => index <= 3;
         when "00111000" => index <= 5;
         when "00111001" => index <= 4;
         when "00111010" => index <= 4;
         when "00111011" => index <= 4;
         when "00111100" => index <= 4;
         when "00111101" => index <= 4;
         when "00111110" => index <= 4;
         when "00111111" => index <= 4;
         when "01000000" => index <= 7;
         when "01000001" => index <= 4;
         when "01000010" => index <= 4;
         when "01000011" => index <= 3;
         when "01000100" => index <= 5;
         when "01000101" => index <= 4;
         when "01000110" => index <= 4;
         when "01000111" => index <= 3;
         when "01001000" => index <= 6;
         when "01001001" => index <= 4;
         when "01001010" => index <= 4;
         when "01001011" => index <= 4;
         when "01001100" => index <= 5;
         when "01001101" => index <= 4;
         when "01001110" => index <= 4;
         when "01001111" => index <= 3;
         when "01010000" => index <= 6;
         when "01010001" => index <= 4;
         when "01010010" => index <= 5;
         when "01010011" => index <= 4;
         when "01010100" => index <= 5;
         when "01010101" => index <= 4;
         when "01010110" => index <= 4;
         when "01010111" => index <= 4;
         when "01011000" => index <= 5;
         when "01011001" => index <= 4;
         when "01011010" => index <= 4;
         when "01011011" => index <= 4;
         when "01011100" => index <= 5;
         when "01011101" => index <= 4;
         when "01011110" => index <= 4;
         when "01011111" => index <= 4;
         when "01100000" => index <= 6;
         when "01100001" => index <= 5;
         when "01100010" => index <= 5;
         when "01100011" => index <= 4;
         when "01100100" => index <= 5;
         when "01100101" => index <= 4;
         when "01100110" => index <= 4;
         when "01100111" => index <= 4;
         when "01101000" => index <= 6;
         when "01101001" => index <= 4;
         when "01101010" => index <= 5;
         when "01101011" => index <= 4;
         when "01101100" => index <= 5;
         when "01101101" => index <= 4;
         when "01101110" => index <= 4;
         when "01101111" => index <= 4;
         when "01110000" => index <= 6;
         when "01110001" => index <= 5;
         when "01110010" => index <= 5;
         when "01110011" => index <= 4;
         when "01110100" => index <= 5;
         when "01110101" => index <= 4;
         when "01110110" => index <= 5;
         when "01110111" => index <= 4;
         when "01111000" => index <= 6;
         when "01111001" => index <= 5;
         when "01111010" => index <= 5;
         when "01111011" => index <= 4;
         when "01111100" => index <= 5;
         when "01111101" => index <= 4;
         when "01111110" => index <= 4;
         when "01111111" => index <= 4;
         when "10000000" => index <= 8;
         when "10000001" => index <= 4;
         when "10000010" => index <= 5;
         when "10000011" => index <= 4;
         when "10000100" => index <= 6;
         when "10000101" => index <= 4;
         when "10000110" => index <= 4;
         when "10000111" => index <= 4;
         when "10001000" => index <= 6;
         when "10001001" => index <= 4;
         when "10001010" => index <= 5;
         when "10001011" => index <= 4;
         when "10001100" => index <= 5;
         when "10001101" => index <= 4;
         when "10001110" => index <= 4;
         when "10001111" => index <= 4;
         when "10010000" => index <= 6;
         when "10010001" => index <= 5;
         when "10010010" => index <= 5;
         when "10010011" => index <= 4;
         when "10010100" => index <= 5;
         when "10010101" => index <= 4;
         when "10010110" => index <= 4;
         when "10010111" => index <= 4;
         when "10011000" => index <= 6;
         when "10011001" => index <= 4;
         when "10011010" => index <= 5;
         when "10011011" => index <= 4;
         when "10011100" => index <= 5;
         when "10011101" => index <= 4;
         when "10011110" => index <= 4;
         when "10011111" => index <= 4;
         when "10100000" => index <= 7;
         when "10100001" => index <= 5;
         when "10100010" => index <= 5;
         when "10100011" => index <= 4;
         when "10100100" => index <= 6;
         when "10100101" => index <= 4;
         when "10100110" => index <= 5;
         when "10100111" => index <= 4;
         when "10101000" => index <= 6;
         when "10101001" => index <= 5;
         when "10101010" => index <= 5;
         when "10101011" => index <= 4;
         when "10101100" => index <= 5;
         when "10101101" => index <= 4;
         when "10101110" => index <= 5;
         when "10101111" => index <= 4;
         when "10110000" => index <= 6;
         when "10110001" => index <= 5;
         when "10110010" => index <= 5;
         when "10110011" => index <= 4;
         when "10110100" => index <= 6;
         when "10110101" => index <= 5;
         when "10110110" => index <= 5;
         when "10110111" => index <= 4;
         when "10111000" => index <= 6;
         when "10111001" => index <= 5;
         when "10111010" => index <= 5;
         when "10111011" => index <= 4;
         when "10111100" => index <= 5;
         when "10111101" => index <= 4;
         when "10111110" => index <= 5;
         when "10111111" => index <= 4;
         when "11000000" => index <= 8;
         when "11000001" => index <= 5;
         when "11000010" => index <= 6;
         when "11000011" => index <= 4;
         when "11000100" => index <= 6;
         when "11000101" => index <= 5;
         when "11000110" => index <= 5;
         when "11000111" => index <= 4;
         when "11001000" => index <= 6;
         when "11001001" => index <= 5;
         when "11001010" => index <= 5;
         when "11001011" => index <= 4;
         when "11001100" => index <= 6;
         when "11001101" => index <= 5;
         when "11001110" => index <= 5;
         when "11001111" => index <= 4;
         when "11010000" => index <= 7;
         when "11010001" => index <= 5;
         when "11010010" => index <= 6;
         when "11010011" => index <= 5;
         when "11010100" => index <= 6;
         when "11010101" => index <= 5;
         when "11010110" => index <= 5;
         when "11010111" => index <= 4;
         when "11011000" => index <= 6;
         when "11011001" => index <= 5;
         when "11011010" => index <= 5;
         when "11011011" => index <= 4;
         when "11011100" => index <= 5;
         when "11011101" => index <= 5;
         when "11011110" => index <= 5;
         when "11011111" => index <= 4;
         when "11100000" => index <= 7;
         when "11100001" => index <= 6;
         when "11100010" => index <= 6;
         when "11100011" => index <= 5;
         when "11100100" => index <= 6;
         when "11100101" => index <= 5;
         when "11100110" => index <= 5;
         when "11100111" => index <= 4;
         when "11101000" => index <= 6;
         when "11101001" => index <= 5;
         when "11101010" => index <= 5;
         when "11101011" => index <= 5;
         when "11101100" => index <= 6;
         when "11101101" => index <= 5;
         when "11101110" => index <= 5;
         when "11101111" => index <= 4;
         when "11110000" => index <= 6;
         when "11110001" => index <= 5;
         when "11110010" => index <= 6;
         when "11110011" => index <= 5;
         when "11110100" => index <= 6;
         when "11110101" => index <= 5;
         when "11110110" => index <= 5;
         when "11110111" => index <= 5;
         when "11111000" => index <= 6;
         when "11111001" => index <= 5;
         when "11111010" => index <= 5;
         when "11111011" => index <= 5;
         when "11111100" => index <= 6;
         when "11111101" => index <= 5;
         when "11111110" => index <= 5;
         when "11111111" => index <= 4;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_9 : if (length = 9) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "000000000" => index <= 0;
         when "000000001" => index <= 1;
         when "000000010" => index <= 2;
         when "000000011" => index <= 2;
         when "000000100" => index <= 3;
         when "000000101" => index <= 2;
         when "000000110" => index <= 2;
         when "000000111" => index <= 2;
         when "000001000" => index <= 4;
         when "000001001" => index <= 2;
         when "000001010" => index <= 3;
         when "000001011" => index <= 2;
         when "000001100" => index <= 4;
         when "000001101" => index <= 3;
         when "000001110" => index <= 3;
         when "000001111" => index <= 2;
         when "000010000" => index <= 5;
         when "000010001" => index <= 3;
         when "000010010" => index <= 4;
         when "000010011" => index <= 3;
         when "000010100" => index <= 4;
         when "000010101" => index <= 3;
         when "000010110" => index <= 3;
         when "000010111" => index <= 3;
         when "000011000" => index <= 4;
         when "000011001" => index <= 3;
         when "000011010" => index <= 4;
         when "000011011" => index <= 3;
         when "000011100" => index <= 4;
         when "000011101" => index <= 3;
         when "000011110" => index <= 4;
         when "000011111" => index <= 3;
         when "000100000" => index <= 6;
         when "000100001" => index <= 4;
         when "000100010" => index <= 4;
         when "000100011" => index <= 3;
         when "000100100" => index <= 4;
         when "000100101" => index <= 3;
         when "000100110" => index <= 4;
         when "000100111" => index <= 3;
         when "000101000" => index <= 5;
         when "000101001" => index <= 4;
         when "000101010" => index <= 4;
         when "000101011" => index <= 3;
         when "000101100" => index <= 4;
         when "000101101" => index <= 4;
         when "000101110" => index <= 4;
         when "000101111" => index <= 3;
         when "000110000" => index <= 6;
         when "000110001" => index <= 4;
         when "000110010" => index <= 4;
         when "000110011" => index <= 4;
         when "000110100" => index <= 5;
         when "000110101" => index <= 4;
         when "000110110" => index <= 4;
         when "000110111" => index <= 3;
         when "000111000" => index <= 5;
         when "000111001" => index <= 4;
         when "000111010" => index <= 4;
         when "000111011" => index <= 4;
         when "000111100" => index <= 4;
         when "000111101" => index <= 4;
         when "000111110" => index <= 4;
         when "000111111" => index <= 4;
         when "001000000" => index <= 7;
         when "001000001" => index <= 4;
         when "001000010" => index <= 4;
         when "001000011" => index <= 3;
         when "001000100" => index <= 5;
         when "001000101" => index <= 4;
         when "001000110" => index <= 4;
         when "001000111" => index <= 3;
         when "001001000" => index <= 6;
         when "001001001" => index <= 4;
         when "001001010" => index <= 4;
         when "001001011" => index <= 4;
         when "001001100" => index <= 5;
         when "001001101" => index <= 4;
         when "001001110" => index <= 4;
         when "001001111" => index <= 3;
         when "001010000" => index <= 6;
         when "001010001" => index <= 4;
         when "001010010" => index <= 5;
         when "001010011" => index <= 4;
         when "001010100" => index <= 5;
         when "001010101" => index <= 4;
         when "001010110" => index <= 4;
         when "001010111" => index <= 4;
         when "001011000" => index <= 5;
         when "001011001" => index <= 4;
         when "001011010" => index <= 4;
         when "001011011" => index <= 4;
         when "001011100" => index <= 5;
         when "001011101" => index <= 4;
         when "001011110" => index <= 4;
         when "001011111" => index <= 4;
         when "001100000" => index <= 6;
         when "001100001" => index <= 5;
         when "001100010" => index <= 5;
         when "001100011" => index <= 4;
         when "001100100" => index <= 5;
         when "001100101" => index <= 4;
         when "001100110" => index <= 4;
         when "001100111" => index <= 4;
         when "001101000" => index <= 6;
         when "001101001" => index <= 4;
         when "001101010" => index <= 5;
         when "001101011" => index <= 4;
         when "001101100" => index <= 5;
         when "001101101" => index <= 4;
         when "001101110" => index <= 4;
         when "001101111" => index <= 4;
         when "001110000" => index <= 6;
         when "001110001" => index <= 5;
         when "001110010" => index <= 5;
         when "001110011" => index <= 4;
         when "001110100" => index <= 5;
         when "001110101" => index <= 4;
         when "001110110" => index <= 5;
         when "001110111" => index <= 4;
         when "001111000" => index <= 6;
         when "001111001" => index <= 5;
         when "001111010" => index <= 5;
         when "001111011" => index <= 4;
         when "001111100" => index <= 5;
         when "001111101" => index <= 4;
         when "001111110" => index <= 4;
         when "001111111" => index <= 4;
         when "010000000" => index <= 8;
         when "010000001" => index <= 4;
         when "010000010" => index <= 5;
         when "010000011" => index <= 4;
         when "010000100" => index <= 6;
         when "010000101" => index <= 4;
         when "010000110" => index <= 4;
         when "010000111" => index <= 4;
         when "010001000" => index <= 6;
         when "010001001" => index <= 4;
         when "010001010" => index <= 5;
         when "010001011" => index <= 4;
         when "010001100" => index <= 5;
         when "010001101" => index <= 4;
         when "010001110" => index <= 4;
         when "010001111" => index <= 4;
         when "010010000" => index <= 6;
         when "010010001" => index <= 5;
         when "010010010" => index <= 5;
         when "010010011" => index <= 4;
         when "010010100" => index <= 5;
         when "010010101" => index <= 4;
         when "010010110" => index <= 4;
         when "010010111" => index <= 4;
         when "010011000" => index <= 6;
         when "010011001" => index <= 4;
         when "010011010" => index <= 5;
         when "010011011" => index <= 4;
         when "010011100" => index <= 5;
         when "010011101" => index <= 4;
         when "010011110" => index <= 4;
         when "010011111" => index <= 4;
         when "010100000" => index <= 7;
         when "010100001" => index <= 5;
         when "010100010" => index <= 5;
         when "010100011" => index <= 4;
         when "010100100" => index <= 6;
         when "010100101" => index <= 4;
         when "010100110" => index <= 5;
         when "010100111" => index <= 4;
         when "010101000" => index <= 6;
         when "010101001" => index <= 5;
         when "010101010" => index <= 5;
         when "010101011" => index <= 4;
         when "010101100" => index <= 5;
         when "010101101" => index <= 4;
         when "010101110" => index <= 5;
         when "010101111" => index <= 4;
         when "010110000" => index <= 6;
         when "010110001" => index <= 5;
         when "010110010" => index <= 5;
         when "010110011" => index <= 4;
         when "010110100" => index <= 6;
         when "010110101" => index <= 5;
         when "010110110" => index <= 5;
         when "010110111" => index <= 4;
         when "010111000" => index <= 6;
         when "010111001" => index <= 5;
         when "010111010" => index <= 5;
         when "010111011" => index <= 4;
         when "010111100" => index <= 5;
         when "010111101" => index <= 4;
         when "010111110" => index <= 5;
         when "010111111" => index <= 4;
         when "011000000" => index <= 8;
         when "011000001" => index <= 5;
         when "011000010" => index <= 6;
         when "011000011" => index <= 4;
         when "011000100" => index <= 6;
         when "011000101" => index <= 5;
         when "011000110" => index <= 5;
         when "011000111" => index <= 4;
         when "011001000" => index <= 6;
         when "011001001" => index <= 5;
         when "011001010" => index <= 5;
         when "011001011" => index <= 4;
         when "011001100" => index <= 6;
         when "011001101" => index <= 5;
         when "011001110" => index <= 5;
         when "011001111" => index <= 4;
         when "011010000" => index <= 7;
         when "011010001" => index <= 5;
         when "011010010" => index <= 6;
         when "011010011" => index <= 5;
         when "011010100" => index <= 6;
         when "011010101" => index <= 5;
         when "011010110" => index <= 5;
         when "011010111" => index <= 4;
         when "011011000" => index <= 6;
         when "011011001" => index <= 5;
         when "011011010" => index <= 5;
         when "011011011" => index <= 4;
         when "011011100" => index <= 5;
         when "011011101" => index <= 5;
         when "011011110" => index <= 5;
         when "011011111" => index <= 4;
         when "011100000" => index <= 7;
         when "011100001" => index <= 6;
         when "011100010" => index <= 6;
         when "011100011" => index <= 5;
         when "011100100" => index <= 6;
         when "011100101" => index <= 5;
         when "011100110" => index <= 5;
         when "011100111" => index <= 4;
         when "011101000" => index <= 6;
         when "011101001" => index <= 5;
         when "011101010" => index <= 5;
         when "011101011" => index <= 5;
         when "011101100" => index <= 6;
         when "011101101" => index <= 5;
         when "011101110" => index <= 5;
         when "011101111" => index <= 4;
         when "011110000" => index <= 6;
         when "011110001" => index <= 5;
         when "011110010" => index <= 6;
         when "011110011" => index <= 5;
         when "011110100" => index <= 6;
         when "011110101" => index <= 5;
         when "011110110" => index <= 5;
         when "011110111" => index <= 5;
         when "011111000" => index <= 6;
         when "011111001" => index <= 5;
         when "011111010" => index <= 5;
         when "011111011" => index <= 5;
         when "011111100" => index <= 6;
         when "011111101" => index <= 5;
         when "011111110" => index <= 5;
         when "011111111" => index <= 4;
         when "100000000" => index <= 9;
         when "100000001" => index <= 5;
         when "100000010" => index <= 6;
         when "100000011" => index <= 4;
         when "100000100" => index <= 6;
         when "100000101" => index <= 4;
         when "100000110" => index <= 5;
         when "100000111" => index <= 4;
         when "100001000" => index <= 6;
         when "100001001" => index <= 5;
         when "100001010" => index <= 5;
         when "100001011" => index <= 4;
         when "100001100" => index <= 5;
         when "100001101" => index <= 4;
         when "100001110" => index <= 4;
         when "100001111" => index <= 4;
         when "100010000" => index <= 7;
         when "100010001" => index <= 5;
         when "100010010" => index <= 5;
         when "100010011" => index <= 4;
         when "100010100" => index <= 6;
         when "100010101" => index <= 4;
         when "100010110" => index <= 5;
         when "100010111" => index <= 4;
         when "100011000" => index <= 6;
         when "100011001" => index <= 5;
         when "100011010" => index <= 5;
         when "100011011" => index <= 4;
         when "100011100" => index <= 5;
         when "100011101" => index <= 4;
         when "100011110" => index <= 5;
         when "100011111" => index <= 4;
         when "100100000" => index <= 8;
         when "100100001" => index <= 5;
         when "100100010" => index <= 6;
         when "100100011" => index <= 4;
         when "100100100" => index <= 6;
         when "100100101" => index <= 5;
         when "100100110" => index <= 5;
         when "100100111" => index <= 4;
         when "100101000" => index <= 6;
         when "100101001" => index <= 5;
         when "100101010" => index <= 5;
         when "100101011" => index <= 4;
         when "100101100" => index <= 6;
         when "100101101" => index <= 5;
         when "100101110" => index <= 5;
         when "100101111" => index <= 4;
         when "100110000" => index <= 7;
         when "100110001" => index <= 5;
         when "100110010" => index <= 6;
         when "100110011" => index <= 5;
         when "100110100" => index <= 6;
         when "100110101" => index <= 5;
         when "100110110" => index <= 5;
         when "100110111" => index <= 4;
         when "100111000" => index <= 6;
         when "100111001" => index <= 5;
         when "100111010" => index <= 5;
         when "100111011" => index <= 4;
         when "100111100" => index <= 5;
         when "100111101" => index <= 5;
         when "100111110" => index <= 5;
         when "100111111" => index <= 4;
         when "101000000" => index <= 8;
         when "101000001" => index <= 6;
         when "101000010" => index <= 6;
         when "101000011" => index <= 5;
         when "101000100" => index <= 6;
         when "101000101" => index <= 5;
         when "101000110" => index <= 5;
         when "101000111" => index <= 4;
         when "101001000" => index <= 7;
         when "101001001" => index <= 5;
         when "101001010" => index <= 6;
         when "101001011" => index <= 5;
         when "101001100" => index <= 6;
         when "101001101" => index <= 5;
         when "101001110" => index <= 5;
         when "101001111" => index <= 4;
         when "101010000" => index <= 7;
         when "101010001" => index <= 6;
         when "101010010" => index <= 6;
         when "101010011" => index <= 5;
         when "101010100" => index <= 6;
         when "101010101" => index <= 5;
         when "101010110" => index <= 5;
         when "101010111" => index <= 4;
         when "101011000" => index <= 6;
         when "101011001" => index <= 5;
         when "101011010" => index <= 5;
         when "101011011" => index <= 5;
         when "101011100" => index <= 6;
         when "101011101" => index <= 5;
         when "101011110" => index <= 5;
         when "101011111" => index <= 4;
         when "101100000" => index <= 7;
         when "101100001" => index <= 6;
         when "101100010" => index <= 6;
         when "101100011" => index <= 5;
         when "101100100" => index <= 6;
         when "101100101" => index <= 5;
         when "101100110" => index <= 5;
         when "101100111" => index <= 5;
         when "101101000" => index <= 6;
         when "101101001" => index <= 5;
         when "101101010" => index <= 6;
         when "101101011" => index <= 5;
         when "101101100" => index <= 6;
         when "101101101" => index <= 5;
         when "101101110" => index <= 5;
         when "101101111" => index <= 5;
         when "101110000" => index <= 7;
         when "101110001" => index <= 6;
         when "101110010" => index <= 6;
         when "101110011" => index <= 5;
         when "101110100" => index <= 6;
         when "101110101" => index <= 5;
         when "101110110" => index <= 5;
         when "101110111" => index <= 5;
         when "101111000" => index <= 6;
         when "101111001" => index <= 5;
         when "101111010" => index <= 6;
         when "101111011" => index <= 5;
         when "101111100" => index <= 6;
         when "101111101" => index <= 5;
         when "101111110" => index <= 5;
         when "101111111" => index <= 5;
         when "110000000" => index <= 8;
         when "110000001" => index <= 6;
         when "110000010" => index <= 6;
         when "110000011" => index <= 5;
         when "110000100" => index <= 7;
         when "110000101" => index <= 5;
         when "110000110" => index <= 6;
         when "110000111" => index <= 5;
         when "110001000" => index <= 7;
         when "110001001" => index <= 6;
         when "110001010" => index <= 6;
         when "110001011" => index <= 5;
         when "110001100" => index <= 6;
         when "110001101" => index <= 5;
         when "110001110" => index <= 5;
         when "110001111" => index <= 4;
         when "110010000" => index <= 7;
         when "110010001" => index <= 6;
         when "110010010" => index <= 6;
         when "110010011" => index <= 5;
         when "110010100" => index <= 6;
         when "110010101" => index <= 5;
         when "110010110" => index <= 5;
         when "110010111" => index <= 5;
         when "110011000" => index <= 6;
         when "110011001" => index <= 5;
         when "110011010" => index <= 6;
         when "110011011" => index <= 5;
         when "110011100" => index <= 6;
         when "110011101" => index <= 5;
         when "110011110" => index <= 5;
         when "110011111" => index <= 5;
         when "110100000" => index <= 8;
         when "110100001" => index <= 6;
         when "110100010" => index <= 6;
         when "110100011" => index <= 5;
         when "110100100" => index <= 6;
         when "110100101" => index <= 5;
         when "110100110" => index <= 6;
         when "110100111" => index <= 5;
         when "110101000" => index <= 7;
         when "110101001" => index <= 6;
         when "110101010" => index <= 6;
         when "110101011" => index <= 5;
         when "110101100" => index <= 6;
         when "110101101" => index <= 5;
         when "110101110" => index <= 5;
         when "110101111" => index <= 5;
         when "110110000" => index <= 7;
         when "110110001" => index <= 6;
         when "110110010" => index <= 6;
         when "110110011" => index <= 5;
         when "110110100" => index <= 6;
         when "110110101" => index <= 5;
         when "110110110" => index <= 6;
         when "110110111" => index <= 5;
         when "110111000" => index <= 6;
         when "110111001" => index <= 6;
         when "110111010" => index <= 6;
         when "110111011" => index <= 5;
         when "110111100" => index <= 6;
         when "110111101" => index <= 5;
         when "110111110" => index <= 5;
         when "110111111" => index <= 5;
         when "111000000" => index <= 8;
         when "111000001" => index <= 6;
         when "111000010" => index <= 6;
         when "111000011" => index <= 5;
         when "111000100" => index <= 7;
         when "111000101" => index <= 6;
         when "111000110" => index <= 6;
         when "111000111" => index <= 5;
         when "111001000" => index <= 7;
         when "111001001" => index <= 6;
         when "111001010" => index <= 6;
         when "111001011" => index <= 5;
         when "111001100" => index <= 6;
         when "111001101" => index <= 5;
         when "111001110" => index <= 6;
         when "111001111" => index <= 5;
         when "111010000" => index <= 7;
         when "111010001" => index <= 6;
         when "111010010" => index <= 6;
         when "111010011" => index <= 5;
         when "111010100" => index <= 6;
         when "111010101" => index <= 6;
         when "111010110" => index <= 6;
         when "111010111" => index <= 5;
         when "111011000" => index <= 7;
         when "111011001" => index <= 6;
         when "111011010" => index <= 6;
         when "111011011" => index <= 5;
         when "111011100" => index <= 6;
         when "111011101" => index <= 5;
         when "111011110" => index <= 5;
         when "111011111" => index <= 5;
         when "111100000" => index <= 8;
         when "111100001" => index <= 6;
         when "111100010" => index <= 6;
         when "111100011" => index <= 6;
         when "111100100" => index <= 7;
         when "111100101" => index <= 6;
         when "111100110" => index <= 6;
         when "111100111" => index <= 5;
         when "111101000" => index <= 7;
         when "111101001" => index <= 6;
         when "111101010" => index <= 6;
         when "111101011" => index <= 5;
         when "111101100" => index <= 6;
         when "111101101" => index <= 5;
         when "111101110" => index <= 6;
         when "111101111" => index <= 5;
         when "111110000" => index <= 7;
         when "111110001" => index <= 6;
         when "111110010" => index <= 6;
         when "111110011" => index <= 5;
         when "111110100" => index <= 6;
         when "111110101" => index <= 6;
         when "111110110" => index <= 6;
         when "111110111" => index <= 5;
         when "111111000" => index <= 6;
         when "111111001" => index <= 6;
         when "111111010" => index <= 6;
         when "111111011" => index <= 5;
         when "111111100" => index <= 6;
         when "111111101" => index <= 5;
         when "111111110" => index <= 6;
         when "111111111" => index <= 5;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_10 : if (length = 10) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "0000000000" => index <= 0;
         when "0000000001" => index <= 1;
         when "0000000010" => index <= 2;
         when "0000000011" => index <= 2;
         when "0000000100" => index <= 3;
         when "0000000101" => index <= 2;
         when "0000000110" => index <= 2;
         when "0000000111" => index <= 2;
         when "0000001000" => index <= 4;
         when "0000001001" => index <= 2;
         when "0000001010" => index <= 3;
         when "0000001011" => index <= 2;
         when "0000001100" => index <= 4;
         when "0000001101" => index <= 3;
         when "0000001110" => index <= 3;
         when "0000001111" => index <= 2;
         when "0000010000" => index <= 5;
         when "0000010001" => index <= 3;
         when "0000010010" => index <= 4;
         when "0000010011" => index <= 3;
         when "0000010100" => index <= 4;
         when "0000010101" => index <= 3;
         when "0000010110" => index <= 3;
         when "0000010111" => index <= 3;
         when "0000011000" => index <= 4;
         when "0000011001" => index <= 3;
         when "0000011010" => index <= 4;
         when "0000011011" => index <= 3;
         when "0000011100" => index <= 4;
         when "0000011101" => index <= 3;
         when "0000011110" => index <= 4;
         when "0000011111" => index <= 3;
         when "0000100000" => index <= 6;
         when "0000100001" => index <= 4;
         when "0000100010" => index <= 4;
         when "0000100011" => index <= 3;
         when "0000100100" => index <= 4;
         when "0000100101" => index <= 3;
         when "0000100110" => index <= 4;
         when "0000100111" => index <= 3;
         when "0000101000" => index <= 5;
         when "0000101001" => index <= 4;
         when "0000101010" => index <= 4;
         when "0000101011" => index <= 3;
         when "0000101100" => index <= 4;
         when "0000101101" => index <= 4;
         when "0000101110" => index <= 4;
         when "0000101111" => index <= 3;
         when "0000110000" => index <= 6;
         when "0000110001" => index <= 4;
         when "0000110010" => index <= 4;
         when "0000110011" => index <= 4;
         when "0000110100" => index <= 5;
         when "0000110101" => index <= 4;
         when "0000110110" => index <= 4;
         when "0000110111" => index <= 3;
         when "0000111000" => index <= 5;
         when "0000111001" => index <= 4;
         when "0000111010" => index <= 4;
         when "0000111011" => index <= 4;
         when "0000111100" => index <= 4;
         when "0000111101" => index <= 4;
         when "0000111110" => index <= 4;
         when "0000111111" => index <= 4;
         when "0001000000" => index <= 7;
         when "0001000001" => index <= 4;
         when "0001000010" => index <= 4;
         when "0001000011" => index <= 3;
         when "0001000100" => index <= 5;
         when "0001000101" => index <= 4;
         when "0001000110" => index <= 4;
         when "0001000111" => index <= 3;
         when "0001001000" => index <= 6;
         when "0001001001" => index <= 4;
         when "0001001010" => index <= 4;
         when "0001001011" => index <= 4;
         when "0001001100" => index <= 5;
         when "0001001101" => index <= 4;
         when "0001001110" => index <= 4;
         when "0001001111" => index <= 3;
         when "0001010000" => index <= 6;
         when "0001010001" => index <= 4;
         when "0001010010" => index <= 5;
         when "0001010011" => index <= 4;
         when "0001010100" => index <= 5;
         when "0001010101" => index <= 4;
         when "0001010110" => index <= 4;
         when "0001010111" => index <= 4;
         when "0001011000" => index <= 5;
         when "0001011001" => index <= 4;
         when "0001011010" => index <= 4;
         when "0001011011" => index <= 4;
         when "0001011100" => index <= 5;
         when "0001011101" => index <= 4;
         when "0001011110" => index <= 4;
         when "0001011111" => index <= 4;
         when "0001100000" => index <= 6;
         when "0001100001" => index <= 5;
         when "0001100010" => index <= 5;
         when "0001100011" => index <= 4;
         when "0001100100" => index <= 5;
         when "0001100101" => index <= 4;
         when "0001100110" => index <= 4;
         when "0001100111" => index <= 4;
         when "0001101000" => index <= 6;
         when "0001101001" => index <= 4;
         when "0001101010" => index <= 5;
         when "0001101011" => index <= 4;
         when "0001101100" => index <= 5;
         when "0001101101" => index <= 4;
         when "0001101110" => index <= 4;
         when "0001101111" => index <= 4;
         when "0001110000" => index <= 6;
         when "0001110001" => index <= 5;
         when "0001110010" => index <= 5;
         when "0001110011" => index <= 4;
         when "0001110100" => index <= 5;
         when "0001110101" => index <= 4;
         when "0001110110" => index <= 5;
         when "0001110111" => index <= 4;
         when "0001111000" => index <= 6;
         when "0001111001" => index <= 5;
         when "0001111010" => index <= 5;
         when "0001111011" => index <= 4;
         when "0001111100" => index <= 5;
         when "0001111101" => index <= 4;
         when "0001111110" => index <= 4;
         when "0001111111" => index <= 4;
         when "0010000000" => index <= 8;
         when "0010000001" => index <= 4;
         when "0010000010" => index <= 5;
         when "0010000011" => index <= 4;
         when "0010000100" => index <= 6;
         when "0010000101" => index <= 4;
         when "0010000110" => index <= 4;
         when "0010000111" => index <= 4;
         when "0010001000" => index <= 6;
         when "0010001001" => index <= 4;
         when "0010001010" => index <= 5;
         when "0010001011" => index <= 4;
         when "0010001100" => index <= 5;
         when "0010001101" => index <= 4;
         when "0010001110" => index <= 4;
         when "0010001111" => index <= 4;
         when "0010010000" => index <= 6;
         when "0010010001" => index <= 5;
         when "0010010010" => index <= 5;
         when "0010010011" => index <= 4;
         when "0010010100" => index <= 5;
         when "0010010101" => index <= 4;
         when "0010010110" => index <= 4;
         when "0010010111" => index <= 4;
         when "0010011000" => index <= 6;
         when "0010011001" => index <= 4;
         when "0010011010" => index <= 5;
         when "0010011011" => index <= 4;
         when "0010011100" => index <= 5;
         when "0010011101" => index <= 4;
         when "0010011110" => index <= 4;
         when "0010011111" => index <= 4;
         when "0010100000" => index <= 7;
         when "0010100001" => index <= 5;
         when "0010100010" => index <= 5;
         when "0010100011" => index <= 4;
         when "0010100100" => index <= 6;
         when "0010100101" => index <= 4;
         when "0010100110" => index <= 5;
         when "0010100111" => index <= 4;
         when "0010101000" => index <= 6;
         when "0010101001" => index <= 5;
         when "0010101010" => index <= 5;
         when "0010101011" => index <= 4;
         when "0010101100" => index <= 5;
         when "0010101101" => index <= 4;
         when "0010101110" => index <= 5;
         when "0010101111" => index <= 4;
         when "0010110000" => index <= 6;
         when "0010110001" => index <= 5;
         when "0010110010" => index <= 5;
         when "0010110011" => index <= 4;
         when "0010110100" => index <= 6;
         when "0010110101" => index <= 5;
         when "0010110110" => index <= 5;
         when "0010110111" => index <= 4;
         when "0010111000" => index <= 6;
         when "0010111001" => index <= 5;
         when "0010111010" => index <= 5;
         when "0010111011" => index <= 4;
         when "0010111100" => index <= 5;
         when "0010111101" => index <= 4;
         when "0010111110" => index <= 5;
         when "0010111111" => index <= 4;
         when "0011000000" => index <= 8;
         when "0011000001" => index <= 5;
         when "0011000010" => index <= 6;
         when "0011000011" => index <= 4;
         when "0011000100" => index <= 6;
         when "0011000101" => index <= 5;
         when "0011000110" => index <= 5;
         when "0011000111" => index <= 4;
         when "0011001000" => index <= 6;
         when "0011001001" => index <= 5;
         when "0011001010" => index <= 5;
         when "0011001011" => index <= 4;
         when "0011001100" => index <= 6;
         when "0011001101" => index <= 5;
         when "0011001110" => index <= 5;
         when "0011001111" => index <= 4;
         when "0011010000" => index <= 7;
         when "0011010001" => index <= 5;
         when "0011010010" => index <= 6;
         when "0011010011" => index <= 5;
         when "0011010100" => index <= 6;
         when "0011010101" => index <= 5;
         when "0011010110" => index <= 5;
         when "0011010111" => index <= 4;
         when "0011011000" => index <= 6;
         when "0011011001" => index <= 5;
         when "0011011010" => index <= 5;
         when "0011011011" => index <= 4;
         when "0011011100" => index <= 5;
         when "0011011101" => index <= 5;
         when "0011011110" => index <= 5;
         when "0011011111" => index <= 4;
         when "0011100000" => index <= 7;
         when "0011100001" => index <= 6;
         when "0011100010" => index <= 6;
         when "0011100011" => index <= 5;
         when "0011100100" => index <= 6;
         when "0011100101" => index <= 5;
         when "0011100110" => index <= 5;
         when "0011100111" => index <= 4;
         when "0011101000" => index <= 6;
         when "0011101001" => index <= 5;
         when "0011101010" => index <= 5;
         when "0011101011" => index <= 5;
         when "0011101100" => index <= 6;
         when "0011101101" => index <= 5;
         when "0011101110" => index <= 5;
         when "0011101111" => index <= 4;
         when "0011110000" => index <= 6;
         when "0011110001" => index <= 5;
         when "0011110010" => index <= 6;
         when "0011110011" => index <= 5;
         when "0011110100" => index <= 6;
         when "0011110101" => index <= 5;
         when "0011110110" => index <= 5;
         when "0011110111" => index <= 5;
         when "0011111000" => index <= 6;
         when "0011111001" => index <= 5;
         when "0011111010" => index <= 5;
         when "0011111011" => index <= 5;
         when "0011111100" => index <= 6;
         when "0011111101" => index <= 5;
         when "0011111110" => index <= 5;
         when "0011111111" => index <= 4;
         when "0100000000" => index <= 9;
         when "0100000001" => index <= 5;
         when "0100000010" => index <= 6;
         when "0100000011" => index <= 4;
         when "0100000100" => index <= 6;
         when "0100000101" => index <= 4;
         when "0100000110" => index <= 5;
         when "0100000111" => index <= 4;
         when "0100001000" => index <= 6;
         when "0100001001" => index <= 5;
         when "0100001010" => index <= 5;
         when "0100001011" => index <= 4;
         when "0100001100" => index <= 5;
         when "0100001101" => index <= 4;
         when "0100001110" => index <= 4;
         when "0100001111" => index <= 4;
         when "0100010000" => index <= 7;
         when "0100010001" => index <= 5;
         when "0100010010" => index <= 5;
         when "0100010011" => index <= 4;
         when "0100010100" => index <= 6;
         when "0100010101" => index <= 4;
         when "0100010110" => index <= 5;
         when "0100010111" => index <= 4;
         when "0100011000" => index <= 6;
         when "0100011001" => index <= 5;
         when "0100011010" => index <= 5;
         when "0100011011" => index <= 4;
         when "0100011100" => index <= 5;
         when "0100011101" => index <= 4;
         when "0100011110" => index <= 5;
         when "0100011111" => index <= 4;
         when "0100100000" => index <= 8;
         when "0100100001" => index <= 5;
         when "0100100010" => index <= 6;
         when "0100100011" => index <= 4;
         when "0100100100" => index <= 6;
         when "0100100101" => index <= 5;
         when "0100100110" => index <= 5;
         when "0100100111" => index <= 4;
         when "0100101000" => index <= 6;
         when "0100101001" => index <= 5;
         when "0100101010" => index <= 5;
         when "0100101011" => index <= 4;
         when "0100101100" => index <= 6;
         when "0100101101" => index <= 5;
         when "0100101110" => index <= 5;
         when "0100101111" => index <= 4;
         when "0100110000" => index <= 7;
         when "0100110001" => index <= 5;
         when "0100110010" => index <= 6;
         when "0100110011" => index <= 5;
         when "0100110100" => index <= 6;
         when "0100110101" => index <= 5;
         when "0100110110" => index <= 5;
         when "0100110111" => index <= 4;
         when "0100111000" => index <= 6;
         when "0100111001" => index <= 5;
         when "0100111010" => index <= 5;
         when "0100111011" => index <= 4;
         when "0100111100" => index <= 5;
         when "0100111101" => index <= 5;
         when "0100111110" => index <= 5;
         when "0100111111" => index <= 4;
         when "0101000000" => index <= 8;
         when "0101000001" => index <= 6;
         when "0101000010" => index <= 6;
         when "0101000011" => index <= 5;
         when "0101000100" => index <= 6;
         when "0101000101" => index <= 5;
         when "0101000110" => index <= 5;
         when "0101000111" => index <= 4;
         when "0101001000" => index <= 7;
         when "0101001001" => index <= 5;
         when "0101001010" => index <= 6;
         when "0101001011" => index <= 5;
         when "0101001100" => index <= 6;
         when "0101001101" => index <= 5;
         when "0101001110" => index <= 5;
         when "0101001111" => index <= 4;
         when "0101010000" => index <= 7;
         when "0101010001" => index <= 6;
         when "0101010010" => index <= 6;
         when "0101010011" => index <= 5;
         when "0101010100" => index <= 6;
         when "0101010101" => index <= 5;
         when "0101010110" => index <= 5;
         when "0101010111" => index <= 4;
         when "0101011000" => index <= 6;
         when "0101011001" => index <= 5;
         when "0101011010" => index <= 5;
         when "0101011011" => index <= 5;
         when "0101011100" => index <= 6;
         when "0101011101" => index <= 5;
         when "0101011110" => index <= 5;
         when "0101011111" => index <= 4;
         when "0101100000" => index <= 7;
         when "0101100001" => index <= 6;
         when "0101100010" => index <= 6;
         when "0101100011" => index <= 5;
         when "0101100100" => index <= 6;
         when "0101100101" => index <= 5;
         when "0101100110" => index <= 5;
         when "0101100111" => index <= 5;
         when "0101101000" => index <= 6;
         when "0101101001" => index <= 5;
         when "0101101010" => index <= 6;
         when "0101101011" => index <= 5;
         when "0101101100" => index <= 6;
         when "0101101101" => index <= 5;
         when "0101101110" => index <= 5;
         when "0101101111" => index <= 5;
         when "0101110000" => index <= 7;
         when "0101110001" => index <= 6;
         when "0101110010" => index <= 6;
         when "0101110011" => index <= 5;
         when "0101110100" => index <= 6;
         when "0101110101" => index <= 5;
         when "0101110110" => index <= 5;
         when "0101110111" => index <= 5;
         when "0101111000" => index <= 6;
         when "0101111001" => index <= 5;
         when "0101111010" => index <= 6;
         when "0101111011" => index <= 5;
         when "0101111100" => index <= 6;
         when "0101111101" => index <= 5;
         when "0101111110" => index <= 5;
         when "0101111111" => index <= 5;
         when "0110000000" => index <= 8;
         when "0110000001" => index <= 6;
         when "0110000010" => index <= 6;
         when "0110000011" => index <= 5;
         when "0110000100" => index <= 7;
         when "0110000101" => index <= 5;
         when "0110000110" => index <= 6;
         when "0110000111" => index <= 5;
         when "0110001000" => index <= 7;
         when "0110001001" => index <= 6;
         when "0110001010" => index <= 6;
         when "0110001011" => index <= 5;
         when "0110001100" => index <= 6;
         when "0110001101" => index <= 5;
         when "0110001110" => index <= 5;
         when "0110001111" => index <= 4;
         when "0110010000" => index <= 7;
         when "0110010001" => index <= 6;
         when "0110010010" => index <= 6;
         when "0110010011" => index <= 5;
         when "0110010100" => index <= 6;
         when "0110010101" => index <= 5;
         when "0110010110" => index <= 5;
         when "0110010111" => index <= 5;
         when "0110011000" => index <= 6;
         when "0110011001" => index <= 5;
         when "0110011010" => index <= 6;
         when "0110011011" => index <= 5;
         when "0110011100" => index <= 6;
         when "0110011101" => index <= 5;
         when "0110011110" => index <= 5;
         when "0110011111" => index <= 5;
         when "0110100000" => index <= 8;
         when "0110100001" => index <= 6;
         when "0110100010" => index <= 6;
         when "0110100011" => index <= 5;
         when "0110100100" => index <= 6;
         when "0110100101" => index <= 5;
         when "0110100110" => index <= 6;
         when "0110100111" => index <= 5;
         when "0110101000" => index <= 7;
         when "0110101001" => index <= 6;
         when "0110101010" => index <= 6;
         when "0110101011" => index <= 5;
         when "0110101100" => index <= 6;
         when "0110101101" => index <= 5;
         when "0110101110" => index <= 5;
         when "0110101111" => index <= 5;
         when "0110110000" => index <= 7;
         when "0110110001" => index <= 6;
         when "0110110010" => index <= 6;
         when "0110110011" => index <= 5;
         when "0110110100" => index <= 6;
         when "0110110101" => index <= 5;
         when "0110110110" => index <= 6;
         when "0110110111" => index <= 5;
         when "0110111000" => index <= 6;
         when "0110111001" => index <= 6;
         when "0110111010" => index <= 6;
         when "0110111011" => index <= 5;
         when "0110111100" => index <= 6;
         when "0110111101" => index <= 5;
         when "0110111110" => index <= 5;
         when "0110111111" => index <= 5;
         when "0111000000" => index <= 8;
         when "0111000001" => index <= 6;
         when "0111000010" => index <= 6;
         when "0111000011" => index <= 5;
         when "0111000100" => index <= 7;
         when "0111000101" => index <= 6;
         when "0111000110" => index <= 6;
         when "0111000111" => index <= 5;
         when "0111001000" => index <= 7;
         when "0111001001" => index <= 6;
         when "0111001010" => index <= 6;
         when "0111001011" => index <= 5;
         when "0111001100" => index <= 6;
         when "0111001101" => index <= 5;
         when "0111001110" => index <= 6;
         when "0111001111" => index <= 5;
         when "0111010000" => index <= 7;
         when "0111010001" => index <= 6;
         when "0111010010" => index <= 6;
         when "0111010011" => index <= 5;
         when "0111010100" => index <= 6;
         when "0111010101" => index <= 6;
         when "0111010110" => index <= 6;
         when "0111010111" => index <= 5;
         when "0111011000" => index <= 7;
         when "0111011001" => index <= 6;
         when "0111011010" => index <= 6;
         when "0111011011" => index <= 5;
         when "0111011100" => index <= 6;
         when "0111011101" => index <= 5;
         when "0111011110" => index <= 5;
         when "0111011111" => index <= 5;
         when "0111100000" => index <= 8;
         when "0111100001" => index <= 6;
         when "0111100010" => index <= 6;
         when "0111100011" => index <= 6;
         when "0111100100" => index <= 7;
         when "0111100101" => index <= 6;
         when "0111100110" => index <= 6;
         when "0111100111" => index <= 5;
         when "0111101000" => index <= 7;
         when "0111101001" => index <= 6;
         when "0111101010" => index <= 6;
         when "0111101011" => index <= 5;
         when "0111101100" => index <= 6;
         when "0111101101" => index <= 5;
         when "0111101110" => index <= 6;
         when "0111101111" => index <= 5;
         when "0111110000" => index <= 7;
         when "0111110001" => index <= 6;
         when "0111110010" => index <= 6;
         when "0111110011" => index <= 5;
         when "0111110100" => index <= 6;
         when "0111110101" => index <= 6;
         when "0111110110" => index <= 6;
         when "0111110111" => index <= 5;
         when "0111111000" => index <= 6;
         when "0111111001" => index <= 6;
         when "0111111010" => index <= 6;
         when "0111111011" => index <= 5;
         when "0111111100" => index <= 6;
         when "0111111101" => index <= 5;
         when "0111111110" => index <= 6;
         when "0111111111" => index <= 5;
         when "1000000000" => index <= 10;
         when "1000000001" => index <= 6;
         when "1000000010" => index <= 6;
         when "1000000011" => index <= 4;
         when "1000000100" => index <= 6;
         when "1000000101" => index <= 5;
         when "1000000110" => index <= 5;
         when "1000000111" => index <= 4;
         when "1000001000" => index <= 7;
         when "1000001001" => index <= 5;
         when "1000001010" => index <= 5;
         when "1000001011" => index <= 4;
         when "1000001100" => index <= 6;
         when "1000001101" => index <= 4;
         when "1000001110" => index <= 5;
         when "1000001111" => index <= 4;
         when "1000010000" => index <= 8;
         when "1000010001" => index <= 5;
         when "1000010010" => index <= 6;
         when "1000010011" => index <= 4;
         when "1000010100" => index <= 6;
         when "1000010101" => index <= 5;
         when "1000010110" => index <= 5;
         when "1000010111" => index <= 4;
         when "1000011000" => index <= 6;
         when "1000011001" => index <= 5;
         when "1000011010" => index <= 5;
         when "1000011011" => index <= 4;
         when "1000011100" => index <= 6;
         when "1000011101" => index <= 5;
         when "1000011110" => index <= 5;
         when "1000011111" => index <= 4;
         when "1000100000" => index <= 8;
         when "1000100001" => index <= 6;
         when "1000100010" => index <= 6;
         when "1000100011" => index <= 5;
         when "1000100100" => index <= 6;
         when "1000100101" => index <= 5;
         when "1000100110" => index <= 5;
         when "1000100111" => index <= 4;
         when "1000101000" => index <= 7;
         when "1000101001" => index <= 5;
         when "1000101010" => index <= 6;
         when "1000101011" => index <= 5;
         when "1000101100" => index <= 6;
         when "1000101101" => index <= 5;
         when "1000101110" => index <= 5;
         when "1000101111" => index <= 4;
         when "1000110000" => index <= 7;
         when "1000110001" => index <= 6;
         when "1000110010" => index <= 6;
         when "1000110011" => index <= 5;
         when "1000110100" => index <= 6;
         when "1000110101" => index <= 5;
         when "1000110110" => index <= 5;
         when "1000110111" => index <= 4;
         when "1000111000" => index <= 6;
         when "1000111001" => index <= 5;
         when "1000111010" => index <= 5;
         when "1000111011" => index <= 5;
         when "1000111100" => index <= 6;
         when "1000111101" => index <= 5;
         when "1000111110" => index <= 5;
         when "1000111111" => index <= 4;
         when "1001000000" => index <= 8;
         when "1001000001" => index <= 6;
         when "1001000010" => index <= 6;
         when "1001000011" => index <= 5;
         when "1001000100" => index <= 7;
         when "1001000101" => index <= 5;
         when "1001000110" => index <= 6;
         when "1001000111" => index <= 5;
         when "1001001000" => index <= 7;
         when "1001001001" => index <= 6;
         when "1001001010" => index <= 6;
         when "1001001011" => index <= 5;
         when "1001001100" => index <= 6;
         when "1001001101" => index <= 5;
         when "1001001110" => index <= 5;
         when "1001001111" => index <= 4;
         when "1001010000" => index <= 7;
         when "1001010001" => index <= 6;
         when "1001010010" => index <= 6;
         when "1001010011" => index <= 5;
         when "1001010100" => index <= 6;
         when "1001010101" => index <= 5;
         when "1001010110" => index <= 5;
         when "1001010111" => index <= 5;
         when "1001011000" => index <= 6;
         when "1001011001" => index <= 5;
         when "1001011010" => index <= 6;
         when "1001011011" => index <= 5;
         when "1001011100" => index <= 6;
         when "1001011101" => index <= 5;
         when "1001011110" => index <= 5;
         when "1001011111" => index <= 5;
         when "1001100000" => index <= 8;
         when "1001100001" => index <= 6;
         when "1001100010" => index <= 6;
         when "1001100011" => index <= 5;
         when "1001100100" => index <= 6;
         when "1001100101" => index <= 5;
         when "1001100110" => index <= 6;
         when "1001100111" => index <= 5;
         when "1001101000" => index <= 7;
         when "1001101001" => index <= 6;
         when "1001101010" => index <= 6;
         when "1001101011" => index <= 5;
         when "1001101100" => index <= 6;
         when "1001101101" => index <= 5;
         when "1001101110" => index <= 5;
         when "1001101111" => index <= 5;
         when "1001110000" => index <= 7;
         when "1001110001" => index <= 6;
         when "1001110010" => index <= 6;
         when "1001110011" => index <= 5;
         when "1001110100" => index <= 6;
         when "1001110101" => index <= 5;
         when "1001110110" => index <= 6;
         when "1001110111" => index <= 5;
         when "1001111000" => index <= 6;
         when "1001111001" => index <= 6;
         when "1001111010" => index <= 6;
         when "1001111011" => index <= 5;
         when "1001111100" => index <= 6;
         when "1001111101" => index <= 5;
         when "1001111110" => index <= 5;
         when "1001111111" => index <= 5;
         when "1010000000" => index <= 9;
         when "1010000001" => index <= 6;
         when "1010000010" => index <= 7;
         when "1010000011" => index <= 5;
         when "1010000100" => index <= 7;
         when "1010000101" => index <= 6;
         when "1010000110" => index <= 6;
         when "1010000111" => index <= 5;
         when "1010001000" => index <= 7;
         when "1010001001" => index <= 6;
         when "1010001010" => index <= 6;
         when "1010001011" => index <= 5;
         when "1010001100" => index <= 6;
         when "1010001101" => index <= 5;
         when "1010001110" => index <= 5;
         when "1010001111" => index <= 5;
         when "1010010000" => index <= 8;
         when "1010010001" => index <= 6;
         when "1010010010" => index <= 6;
         when "1010010011" => index <= 5;
         when "1010010100" => index <= 6;
         when "1010010101" => index <= 5;
         when "1010010110" => index <= 6;
         when "1010010111" => index <= 5;
         when "1010011000" => index <= 7;
         when "1010011001" => index <= 6;
         when "1010011010" => index <= 6;
         when "1010011011" => index <= 5;
         when "1010011100" => index <= 6;
         when "1010011101" => index <= 5;
         when "1010011110" => index <= 5;
         when "1010011111" => index <= 5;
         when "1010100000" => index <= 8;
         when "1010100001" => index <= 6;
         when "1010100010" => index <= 6;
         when "1010100011" => index <= 5;
         when "1010100100" => index <= 7;
         when "1010100101" => index <= 6;
         when "1010100110" => index <= 6;
         when "1010100111" => index <= 5;
         when "1010101000" => index <= 7;
         when "1010101001" => index <= 6;
         when "1010101010" => index <= 6;
         when "1010101011" => index <= 5;
         when "1010101100" => index <= 6;
         when "1010101101" => index <= 5;
         when "1010101110" => index <= 6;
         when "1010101111" => index <= 5;
         when "1010110000" => index <= 7;
         when "1010110001" => index <= 6;
         when "1010110010" => index <= 6;
         when "1010110011" => index <= 5;
         when "1010110100" => index <= 6;
         when "1010110101" => index <= 6;
         when "1010110110" => index <= 6;
         when "1010110111" => index <= 5;
         when "1010111000" => index <= 7;
         when "1010111001" => index <= 6;
         when "1010111010" => index <= 6;
         when "1010111011" => index <= 5;
         when "1010111100" => index <= 6;
         when "1010111101" => index <= 5;
         when "1010111110" => index <= 5;
         when "1010111111" => index <= 5;
         when "1011000000" => index <= 8;
         when "1011000001" => index <= 6;
         when "1011000010" => index <= 7;
         when "1011000011" => index <= 6;
         when "1011000100" => index <= 7;
         when "1011000101" => index <= 6;
         when "1011000110" => index <= 6;
         when "1011000111" => index <= 5;
         when "1011001000" => index <= 7;
         when "1011001001" => index <= 6;
         when "1011001010" => index <= 6;
         when "1011001011" => index <= 5;
         when "1011001100" => index <= 6;
         when "1011001101" => index <= 6;
         when "1011001110" => index <= 6;
         when "1011001111" => index <= 5;
         when "1011010000" => index <= 8;
         when "1011010001" => index <= 6;
         when "1011010010" => index <= 6;
         when "1011010011" => index <= 6;
         when "1011010100" => index <= 7;
         when "1011010101" => index <= 6;
         when "1011010110" => index <= 6;
         when "1011010111" => index <= 5;
         when "1011011000" => index <= 7;
         when "1011011001" => index <= 6;
         when "1011011010" => index <= 6;
         when "1011011011" => index <= 5;
         when "1011011100" => index <= 6;
         when "1011011101" => index <= 5;
         when "1011011110" => index <= 6;
         when "1011011111" => index <= 5;
         when "1011100000" => index <= 8;
         when "1011100001" => index <= 6;
         when "1011100010" => index <= 7;
         when "1011100011" => index <= 6;
         when "1011100100" => index <= 7;
         when "1011100101" => index <= 6;
         when "1011100110" => index <= 6;
         when "1011100111" => index <= 5;
         when "1011101000" => index <= 7;
         when "1011101001" => index <= 6;
         when "1011101010" => index <= 6;
         when "1011101011" => index <= 5;
         when "1011101100" => index <= 6;
         when "1011101101" => index <= 6;
         when "1011101110" => index <= 6;
         when "1011101111" => index <= 5;
         when "1011110000" => index <= 7;
         when "1011110001" => index <= 6;
         when "1011110010" => index <= 6;
         when "1011110011" => index <= 6;
         when "1011110100" => index <= 6;
         when "1011110101" => index <= 6;
         when "1011110110" => index <= 6;
         when "1011110111" => index <= 5;
         when "1011111000" => index <= 7;
         when "1011111001" => index <= 6;
         when "1011111010" => index <= 6;
         when "1011111011" => index <= 5;
         when "1011111100" => index <= 6;
         when "1011111101" => index <= 6;
         when "1011111110" => index <= 6;
         when "1011111111" => index <= 5;
         when "1100000000" => index <= 10;
         when "1100000001" => index <= 7;
         when "1100000010" => index <= 7;
         when "1100000011" => index <= 6;
         when "1100000100" => index <= 7;
         when "1100000101" => index <= 6;
         when "1100000110" => index <= 6;
         when "1100000111" => index <= 5;
         when "1100001000" => index <= 8;
         when "1100001001" => index <= 6;
         when "1100001010" => index <= 6;
         when "1100001011" => index <= 5;
         when "1100001100" => index <= 6;
         when "1100001101" => index <= 5;
         when "1100001110" => index <= 6;
         when "1100001111" => index <= 5;
         when "1100010000" => index <= 8;
         when "1100010001" => index <= 6;
         when "1100010010" => index <= 6;
         when "1100010011" => index <= 5;
         when "1100010100" => index <= 7;
         when "1100010101" => index <= 6;
         when "1100010110" => index <= 6;
         when "1100010111" => index <= 5;
         when "1100011000" => index <= 7;
         when "1100011001" => index <= 6;
         when "1100011010" => index <= 6;
         when "1100011011" => index <= 5;
         when "1100011100" => index <= 6;
         when "1100011101" => index <= 5;
         when "1100011110" => index <= 6;
         when "1100011111" => index <= 5;
         when "1100100000" => index <= 8;
         when "1100100001" => index <= 6;
         when "1100100010" => index <= 7;
         when "1100100011" => index <= 6;
         when "1100100100" => index <= 7;
         when "1100100101" => index <= 6;
         when "1100100110" => index <= 6;
         when "1100100111" => index <= 5;
         when "1100101000" => index <= 7;
         when "1100101001" => index <= 6;
         when "1100101010" => index <= 6;
         when "1100101011" => index <= 5;
         when "1100101100" => index <= 6;
         when "1100101101" => index <= 6;
         when "1100101110" => index <= 6;
         when "1100101111" => index <= 5;
         when "1100110000" => index <= 8;
         when "1100110001" => index <= 6;
         when "1100110010" => index <= 6;
         when "1100110011" => index <= 6;
         when "1100110100" => index <= 7;
         when "1100110101" => index <= 6;
         when "1100110110" => index <= 6;
         when "1100110111" => index <= 5;
         when "1100111000" => index <= 7;
         when "1100111001" => index <= 6;
         when "1100111010" => index <= 6;
         when "1100111011" => index <= 5;
         when "1100111100" => index <= 6;
         when "1100111101" => index <= 5;
         when "1100111110" => index <= 6;
         when "1100111111" => index <= 5;
         when "1101000000" => index <= 9;
         when "1101000001" => index <= 7;
         when "1101000010" => index <= 7;
         when "1101000011" => index <= 6;
         when "1101000100" => index <= 7;
         when "1101000101" => index <= 6;
         when "1101000110" => index <= 6;
         when "1101000111" => index <= 5;
         when "1101001000" => index <= 8;
         when "1101001001" => index <= 6;
         when "1101001010" => index <= 6;
         when "1101001011" => index <= 6;
         when "1101001100" => index <= 7;
         when "1101001101" => index <= 6;
         when "1101001110" => index <= 6;
         when "1101001111" => index <= 5;
         when "1101010000" => index <= 8;
         when "1101010001" => index <= 6;
         when "1101010010" => index <= 7;
         when "1101010011" => index <= 6;
         when "1101010100" => index <= 7;
         when "1101010101" => index <= 6;
         when "1101010110" => index <= 6;
         when "1101010111" => index <= 5;
         when "1101011000" => index <= 7;
         when "1101011001" => index <= 6;
         when "1101011010" => index <= 6;
         when "1101011011" => index <= 5;
         when "1101011100" => index <= 6;
         when "1101011101" => index <= 6;
         when "1101011110" => index <= 6;
         when "1101011111" => index <= 5;
         when "1101100000" => index <= 8;
         when "1101100001" => index <= 7;
         when "1101100010" => index <= 7;
         when "1101100011" => index <= 6;
         when "1101100100" => index <= 7;
         when "1101100101" => index <= 6;
         when "1101100110" => index <= 6;
         when "1101100111" => index <= 5;
         when "1101101000" => index <= 7;
         when "1101101001" => index <= 6;
         when "1101101010" => index <= 6;
         when "1101101011" => index <= 6;
         when "1101101100" => index <= 6;
         when "1101101101" => index <= 6;
         when "1101101110" => index <= 6;
         when "1101101111" => index <= 5;
         when "1101110000" => index <= 7;
         when "1101110001" => index <= 6;
         when "1101110010" => index <= 6;
         when "1101110011" => index <= 6;
         when "1101110100" => index <= 7;
         when "1101110101" => index <= 6;
         when "1101110110" => index <= 6;
         when "1101110111" => index <= 5;
         when "1101111000" => index <= 7;
         when "1101111001" => index <= 6;
         when "1101111010" => index <= 6;
         when "1101111011" => index <= 6;
         when "1101111100" => index <= 6;
         when "1101111101" => index <= 6;
         when "1101111110" => index <= 6;
         when "1101111111" => index <= 5;
         when "1110000000" => index <= 9;
         when "1110000001" => index <= 7;
         when "1110000010" => index <= 7;
         when "1110000011" => index <= 6;
         when "1110000100" => index <= 8;
         when "1110000101" => index <= 6;
         when "1110000110" => index <= 6;
         when "1110000111" => index <= 6;
         when "1110001000" => index <= 8;
         when "1110001001" => index <= 6;
         when "1110001010" => index <= 7;
         when "1110001011" => index <= 6;
         when "1110001100" => index <= 7;
         when "1110001101" => index <= 6;
         when "1110001110" => index <= 6;
         when "1110001111" => index <= 5;
         when "1110010000" => index <= 8;
         when "1110010001" => index <= 7;
         when "1110010010" => index <= 7;
         when "1110010011" => index <= 6;
         when "1110010100" => index <= 7;
         when "1110010101" => index <= 6;
         when "1110010110" => index <= 6;
         when "1110010111" => index <= 5;
         when "1110011000" => index <= 7;
         when "1110011001" => index <= 6;
         when "1110011010" => index <= 6;
         when "1110011011" => index <= 6;
         when "1110011100" => index <= 6;
         when "1110011101" => index <= 6;
         when "1110011110" => index <= 6;
         when "1110011111" => index <= 5;
         when "1110100000" => index <= 8;
         when "1110100001" => index <= 7;
         when "1110100010" => index <= 7;
         when "1110100011" => index <= 6;
         when "1110100100" => index <= 7;
         when "1110100101" => index <= 6;
         when "1110100110" => index <= 6;
         when "1110100111" => index <= 6;
         when "1110101000" => index <= 7;
         when "1110101001" => index <= 6;
         when "1110101010" => index <= 6;
         when "1110101011" => index <= 6;
         when "1110101100" => index <= 7;
         when "1110101101" => index <= 6;
         when "1110101110" => index <= 6;
         when "1110101111" => index <= 5;
         when "1110110000" => index <= 8;
         when "1110110001" => index <= 6;
         when "1110110010" => index <= 7;
         when "1110110011" => index <= 6;
         when "1110110100" => index <= 7;
         when "1110110101" => index <= 6;
         when "1110110110" => index <= 6;
         when "1110110111" => index <= 6;
         when "1110111000" => index <= 7;
         when "1110111001" => index <= 6;
         when "1110111010" => index <= 6;
         when "1110111011" => index <= 6;
         when "1110111100" => index <= 6;
         when "1110111101" => index <= 6;
         when "1110111110" => index <= 6;
         when "1110111111" => index <= 5;
         when "1111000000" => index <= 8;
         when "1111000001" => index <= 7;
         when "1111000010" => index <= 7;
         when "1111000011" => index <= 6;
         when "1111000100" => index <= 7;
         when "1111000101" => index <= 6;
         when "1111000110" => index <= 6;
         when "1111000111" => index <= 6;
         when "1111001000" => index <= 8;
         when "1111001001" => index <= 6;
         when "1111001010" => index <= 7;
         when "1111001011" => index <= 6;
         when "1111001100" => index <= 7;
         when "1111001101" => index <= 6;
         when "1111001110" => index <= 6;
         when "1111001111" => index <= 6;
         when "1111010000" => index <= 8;
         when "1111010001" => index <= 7;
         when "1111010010" => index <= 7;
         when "1111010011" => index <= 6;
         when "1111010100" => index <= 7;
         when "1111010101" => index <= 6;
         when "1111010110" => index <= 6;
         when "1111010111" => index <= 6;
         when "1111011000" => index <= 7;
         when "1111011001" => index <= 6;
         when "1111011010" => index <= 6;
         when "1111011011" => index <= 6;
         when "1111011100" => index <= 7;
         when "1111011101" => index <= 6;
         when "1111011110" => index <= 6;
         when "1111011111" => index <= 5;
         when "1111100000" => index <= 8;
         when "1111100001" => index <= 7;
         when "1111100010" => index <= 7;
         when "1111100011" => index <= 6;
         when "1111100100" => index <= 7;
         when "1111100101" => index <= 6;
         when "1111100110" => index <= 6;
         when "1111100111" => index <= 6;
         when "1111101000" => index <= 7;
         when "1111101001" => index <= 6;
         when "1111101010" => index <= 7;
         when "1111101011" => index <= 6;
         when "1111101100" => index <= 7;
         when "1111101101" => index <= 6;
         when "1111101110" => index <= 6;
         when "1111101111" => index <= 6;
         when "1111110000" => index <= 8;
         when "1111110001" => index <= 7;
         when "1111110010" => index <= 7;
         when "1111110011" => index <= 6;
         when "1111110100" => index <= 7;
         when "1111110101" => index <= 6;
         when "1111110110" => index <= 6;
         when "1111110111" => index <= 6;
         when "1111111000" => index <= 7;
         when "1111111001" => index <= 6;
         when "1111111010" => index <= 6;
         when "1111111011" => index <= 6;
         when "1111111100" => index <= 6;
         when "1111111101" => index <= 6;
         when "1111111110" => index <= 6;
         when "1111111111" => index <= 6;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_11 : if (length = 11) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "00000000000" => index <= 0;
         when "00000000001" => index <= 1;
         when "00000000010" => index <= 2;
         when "00000000011" => index <= 2;
         when "00000000100" => index <= 3;
         when "00000000101" => index <= 2;
         when "00000000110" => index <= 2;
         when "00000000111" => index <= 2;
         when "00000001000" => index <= 4;
         when "00000001001" => index <= 2;
         when "00000001010" => index <= 3;
         when "00000001011" => index <= 2;
         when "00000001100" => index <= 4;
         when "00000001101" => index <= 3;
         when "00000001110" => index <= 3;
         when "00000001111" => index <= 2;
         when "00000010000" => index <= 5;
         when "00000010001" => index <= 3;
         when "00000010010" => index <= 4;
         when "00000010011" => index <= 3;
         when "00000010100" => index <= 4;
         when "00000010101" => index <= 3;
         when "00000010110" => index <= 3;
         when "00000010111" => index <= 3;
         when "00000011000" => index <= 4;
         when "00000011001" => index <= 3;
         when "00000011010" => index <= 4;
         when "00000011011" => index <= 3;
         when "00000011100" => index <= 4;
         when "00000011101" => index <= 3;
         when "00000011110" => index <= 4;
         when "00000011111" => index <= 3;
         when "00000100000" => index <= 6;
         when "00000100001" => index <= 4;
         when "00000100010" => index <= 4;
         when "00000100011" => index <= 3;
         when "00000100100" => index <= 4;
         when "00000100101" => index <= 3;
         when "00000100110" => index <= 4;
         when "00000100111" => index <= 3;
         when "00000101000" => index <= 5;
         when "00000101001" => index <= 4;
         when "00000101010" => index <= 4;
         when "00000101011" => index <= 3;
         when "00000101100" => index <= 4;
         when "00000101101" => index <= 4;
         when "00000101110" => index <= 4;
         when "00000101111" => index <= 3;
         when "00000110000" => index <= 6;
         when "00000110001" => index <= 4;
         when "00000110010" => index <= 4;
         when "00000110011" => index <= 4;
         when "00000110100" => index <= 5;
         when "00000110101" => index <= 4;
         when "00000110110" => index <= 4;
         when "00000110111" => index <= 3;
         when "00000111000" => index <= 5;
         when "00000111001" => index <= 4;
         when "00000111010" => index <= 4;
         when "00000111011" => index <= 4;
         when "00000111100" => index <= 4;
         when "00000111101" => index <= 4;
         when "00000111110" => index <= 4;
         when "00000111111" => index <= 4;
         when "00001000000" => index <= 7;
         when "00001000001" => index <= 4;
         when "00001000010" => index <= 4;
         when "00001000011" => index <= 3;
         when "00001000100" => index <= 5;
         when "00001000101" => index <= 4;
         when "00001000110" => index <= 4;
         when "00001000111" => index <= 3;
         when "00001001000" => index <= 6;
         when "00001001001" => index <= 4;
         when "00001001010" => index <= 4;
         when "00001001011" => index <= 4;
         when "00001001100" => index <= 5;
         when "00001001101" => index <= 4;
         when "00001001110" => index <= 4;
         when "00001001111" => index <= 3;
         when "00001010000" => index <= 6;
         when "00001010001" => index <= 4;
         when "00001010010" => index <= 5;
         when "00001010011" => index <= 4;
         when "00001010100" => index <= 5;
         when "00001010101" => index <= 4;
         when "00001010110" => index <= 4;
         when "00001010111" => index <= 4;
         when "00001011000" => index <= 5;
         when "00001011001" => index <= 4;
         when "00001011010" => index <= 4;
         when "00001011011" => index <= 4;
         when "00001011100" => index <= 5;
         when "00001011101" => index <= 4;
         when "00001011110" => index <= 4;
         when "00001011111" => index <= 4;
         when "00001100000" => index <= 6;
         when "00001100001" => index <= 5;
         when "00001100010" => index <= 5;
         when "00001100011" => index <= 4;
         when "00001100100" => index <= 5;
         when "00001100101" => index <= 4;
         when "00001100110" => index <= 4;
         when "00001100111" => index <= 4;
         when "00001101000" => index <= 6;
         when "00001101001" => index <= 4;
         when "00001101010" => index <= 5;
         when "00001101011" => index <= 4;
         when "00001101100" => index <= 5;
         when "00001101101" => index <= 4;
         when "00001101110" => index <= 4;
         when "00001101111" => index <= 4;
         when "00001110000" => index <= 6;
         when "00001110001" => index <= 5;
         when "00001110010" => index <= 5;
         when "00001110011" => index <= 4;
         when "00001110100" => index <= 5;
         when "00001110101" => index <= 4;
         when "00001110110" => index <= 5;
         when "00001110111" => index <= 4;
         when "00001111000" => index <= 6;
         when "00001111001" => index <= 5;
         when "00001111010" => index <= 5;
         when "00001111011" => index <= 4;
         when "00001111100" => index <= 5;
         when "00001111101" => index <= 4;
         when "00001111110" => index <= 4;
         when "00001111111" => index <= 4;
         when "00010000000" => index <= 8;
         when "00010000001" => index <= 4;
         when "00010000010" => index <= 5;
         when "00010000011" => index <= 4;
         when "00010000100" => index <= 6;
         when "00010000101" => index <= 4;
         when "00010000110" => index <= 4;
         when "00010000111" => index <= 4;
         when "00010001000" => index <= 6;
         when "00010001001" => index <= 4;
         when "00010001010" => index <= 5;
         when "00010001011" => index <= 4;
         when "00010001100" => index <= 5;
         when "00010001101" => index <= 4;
         when "00010001110" => index <= 4;
         when "00010001111" => index <= 4;
         when "00010010000" => index <= 6;
         when "00010010001" => index <= 5;
         when "00010010010" => index <= 5;
         when "00010010011" => index <= 4;
         when "00010010100" => index <= 5;
         when "00010010101" => index <= 4;
         when "00010010110" => index <= 4;
         when "00010010111" => index <= 4;
         when "00010011000" => index <= 6;
         when "00010011001" => index <= 4;
         when "00010011010" => index <= 5;
         when "00010011011" => index <= 4;
         when "00010011100" => index <= 5;
         when "00010011101" => index <= 4;
         when "00010011110" => index <= 4;
         when "00010011111" => index <= 4;
         when "00010100000" => index <= 7;
         when "00010100001" => index <= 5;
         when "00010100010" => index <= 5;
         when "00010100011" => index <= 4;
         when "00010100100" => index <= 6;
         when "00010100101" => index <= 4;
         when "00010100110" => index <= 5;
         when "00010100111" => index <= 4;
         when "00010101000" => index <= 6;
         when "00010101001" => index <= 5;
         when "00010101010" => index <= 5;
         when "00010101011" => index <= 4;
         when "00010101100" => index <= 5;
         when "00010101101" => index <= 4;
         when "00010101110" => index <= 5;
         when "00010101111" => index <= 4;
         when "00010110000" => index <= 6;
         when "00010110001" => index <= 5;
         when "00010110010" => index <= 5;
         when "00010110011" => index <= 4;
         when "00010110100" => index <= 6;
         when "00010110101" => index <= 5;
         when "00010110110" => index <= 5;
         when "00010110111" => index <= 4;
         when "00010111000" => index <= 6;
         when "00010111001" => index <= 5;
         when "00010111010" => index <= 5;
         when "00010111011" => index <= 4;
         when "00010111100" => index <= 5;
         when "00010111101" => index <= 4;
         when "00010111110" => index <= 5;
         when "00010111111" => index <= 4;
         when "00011000000" => index <= 8;
         when "00011000001" => index <= 5;
         when "00011000010" => index <= 6;
         when "00011000011" => index <= 4;
         when "00011000100" => index <= 6;
         when "00011000101" => index <= 5;
         when "00011000110" => index <= 5;
         when "00011000111" => index <= 4;
         when "00011001000" => index <= 6;
         when "00011001001" => index <= 5;
         when "00011001010" => index <= 5;
         when "00011001011" => index <= 4;
         when "00011001100" => index <= 6;
         when "00011001101" => index <= 5;
         when "00011001110" => index <= 5;
         when "00011001111" => index <= 4;
         when "00011010000" => index <= 7;
         when "00011010001" => index <= 5;
         when "00011010010" => index <= 6;
         when "00011010011" => index <= 5;
         when "00011010100" => index <= 6;
         when "00011010101" => index <= 5;
         when "00011010110" => index <= 5;
         when "00011010111" => index <= 4;
         when "00011011000" => index <= 6;
         when "00011011001" => index <= 5;
         when "00011011010" => index <= 5;
         when "00011011011" => index <= 4;
         when "00011011100" => index <= 5;
         when "00011011101" => index <= 5;
         when "00011011110" => index <= 5;
         when "00011011111" => index <= 4;
         when "00011100000" => index <= 7;
         when "00011100001" => index <= 6;
         when "00011100010" => index <= 6;
         when "00011100011" => index <= 5;
         when "00011100100" => index <= 6;
         when "00011100101" => index <= 5;
         when "00011100110" => index <= 5;
         when "00011100111" => index <= 4;
         when "00011101000" => index <= 6;
         when "00011101001" => index <= 5;
         when "00011101010" => index <= 5;
         when "00011101011" => index <= 5;
         when "00011101100" => index <= 6;
         when "00011101101" => index <= 5;
         when "00011101110" => index <= 5;
         when "00011101111" => index <= 4;
         when "00011110000" => index <= 6;
         when "00011110001" => index <= 5;
         when "00011110010" => index <= 6;
         when "00011110011" => index <= 5;
         when "00011110100" => index <= 6;
         when "00011110101" => index <= 5;
         when "00011110110" => index <= 5;
         when "00011110111" => index <= 5;
         when "00011111000" => index <= 6;
         when "00011111001" => index <= 5;
         when "00011111010" => index <= 5;
         when "00011111011" => index <= 5;
         when "00011111100" => index <= 6;
         when "00011111101" => index <= 5;
         when "00011111110" => index <= 5;
         when "00011111111" => index <= 4;
         when "00100000000" => index <= 9;
         when "00100000001" => index <= 5;
         when "00100000010" => index <= 6;
         when "00100000011" => index <= 4;
         when "00100000100" => index <= 6;
         when "00100000101" => index <= 4;
         when "00100000110" => index <= 5;
         when "00100000111" => index <= 4;
         when "00100001000" => index <= 6;
         when "00100001001" => index <= 5;
         when "00100001010" => index <= 5;
         when "00100001011" => index <= 4;
         when "00100001100" => index <= 5;
         when "00100001101" => index <= 4;
         when "00100001110" => index <= 4;
         when "00100001111" => index <= 4;
         when "00100010000" => index <= 7;
         when "00100010001" => index <= 5;
         when "00100010010" => index <= 5;
         when "00100010011" => index <= 4;
         when "00100010100" => index <= 6;
         when "00100010101" => index <= 4;
         when "00100010110" => index <= 5;
         when "00100010111" => index <= 4;
         when "00100011000" => index <= 6;
         when "00100011001" => index <= 5;
         when "00100011010" => index <= 5;
         when "00100011011" => index <= 4;
         when "00100011100" => index <= 5;
         when "00100011101" => index <= 4;
         when "00100011110" => index <= 5;
         when "00100011111" => index <= 4;
         when "00100100000" => index <= 8;
         when "00100100001" => index <= 5;
         when "00100100010" => index <= 6;
         when "00100100011" => index <= 4;
         when "00100100100" => index <= 6;
         when "00100100101" => index <= 5;
         when "00100100110" => index <= 5;
         when "00100100111" => index <= 4;
         when "00100101000" => index <= 6;
         when "00100101001" => index <= 5;
         when "00100101010" => index <= 5;
         when "00100101011" => index <= 4;
         when "00100101100" => index <= 6;
         when "00100101101" => index <= 5;
         when "00100101110" => index <= 5;
         when "00100101111" => index <= 4;
         when "00100110000" => index <= 7;
         when "00100110001" => index <= 5;
         when "00100110010" => index <= 6;
         when "00100110011" => index <= 5;
         when "00100110100" => index <= 6;
         when "00100110101" => index <= 5;
         when "00100110110" => index <= 5;
         when "00100110111" => index <= 4;
         when "00100111000" => index <= 6;
         when "00100111001" => index <= 5;
         when "00100111010" => index <= 5;
         when "00100111011" => index <= 4;
         when "00100111100" => index <= 5;
         when "00100111101" => index <= 5;
         when "00100111110" => index <= 5;
         when "00100111111" => index <= 4;
         when "00101000000" => index <= 8;
         when "00101000001" => index <= 6;
         when "00101000010" => index <= 6;
         when "00101000011" => index <= 5;
         when "00101000100" => index <= 6;
         when "00101000101" => index <= 5;
         when "00101000110" => index <= 5;
         when "00101000111" => index <= 4;
         when "00101001000" => index <= 7;
         when "00101001001" => index <= 5;
         when "00101001010" => index <= 6;
         when "00101001011" => index <= 5;
         when "00101001100" => index <= 6;
         when "00101001101" => index <= 5;
         when "00101001110" => index <= 5;
         when "00101001111" => index <= 4;
         when "00101010000" => index <= 7;
         when "00101010001" => index <= 6;
         when "00101010010" => index <= 6;
         when "00101010011" => index <= 5;
         when "00101010100" => index <= 6;
         when "00101010101" => index <= 5;
         when "00101010110" => index <= 5;
         when "00101010111" => index <= 4;
         when "00101011000" => index <= 6;
         when "00101011001" => index <= 5;
         when "00101011010" => index <= 5;
         when "00101011011" => index <= 5;
         when "00101011100" => index <= 6;
         when "00101011101" => index <= 5;
         when "00101011110" => index <= 5;
         when "00101011111" => index <= 4;
         when "00101100000" => index <= 7;
         when "00101100001" => index <= 6;
         when "00101100010" => index <= 6;
         when "00101100011" => index <= 5;
         when "00101100100" => index <= 6;
         when "00101100101" => index <= 5;
         when "00101100110" => index <= 5;
         when "00101100111" => index <= 5;
         when "00101101000" => index <= 6;
         when "00101101001" => index <= 5;
         when "00101101010" => index <= 6;
         when "00101101011" => index <= 5;
         when "00101101100" => index <= 6;
         when "00101101101" => index <= 5;
         when "00101101110" => index <= 5;
         when "00101101111" => index <= 5;
         when "00101110000" => index <= 7;
         when "00101110001" => index <= 6;
         when "00101110010" => index <= 6;
         when "00101110011" => index <= 5;
         when "00101110100" => index <= 6;
         when "00101110101" => index <= 5;
         when "00101110110" => index <= 5;
         when "00101110111" => index <= 5;
         when "00101111000" => index <= 6;
         when "00101111001" => index <= 5;
         when "00101111010" => index <= 6;
         when "00101111011" => index <= 5;
         when "00101111100" => index <= 6;
         when "00101111101" => index <= 5;
         when "00101111110" => index <= 5;
         when "00101111111" => index <= 5;
         when "00110000000" => index <= 8;
         when "00110000001" => index <= 6;
         when "00110000010" => index <= 6;
         when "00110000011" => index <= 5;
         when "00110000100" => index <= 7;
         when "00110000101" => index <= 5;
         when "00110000110" => index <= 6;
         when "00110000111" => index <= 5;
         when "00110001000" => index <= 7;
         when "00110001001" => index <= 6;
         when "00110001010" => index <= 6;
         when "00110001011" => index <= 5;
         when "00110001100" => index <= 6;
         when "00110001101" => index <= 5;
         when "00110001110" => index <= 5;
         when "00110001111" => index <= 4;
         when "00110010000" => index <= 7;
         when "00110010001" => index <= 6;
         when "00110010010" => index <= 6;
         when "00110010011" => index <= 5;
         when "00110010100" => index <= 6;
         when "00110010101" => index <= 5;
         when "00110010110" => index <= 5;
         when "00110010111" => index <= 5;
         when "00110011000" => index <= 6;
         when "00110011001" => index <= 5;
         when "00110011010" => index <= 6;
         when "00110011011" => index <= 5;
         when "00110011100" => index <= 6;
         when "00110011101" => index <= 5;
         when "00110011110" => index <= 5;
         when "00110011111" => index <= 5;
         when "00110100000" => index <= 8;
         when "00110100001" => index <= 6;
         when "00110100010" => index <= 6;
         when "00110100011" => index <= 5;
         when "00110100100" => index <= 6;
         when "00110100101" => index <= 5;
         when "00110100110" => index <= 6;
         when "00110100111" => index <= 5;
         when "00110101000" => index <= 7;
         when "00110101001" => index <= 6;
         when "00110101010" => index <= 6;
         when "00110101011" => index <= 5;
         when "00110101100" => index <= 6;
         when "00110101101" => index <= 5;
         when "00110101110" => index <= 5;
         when "00110101111" => index <= 5;
         when "00110110000" => index <= 7;
         when "00110110001" => index <= 6;
         when "00110110010" => index <= 6;
         when "00110110011" => index <= 5;
         when "00110110100" => index <= 6;
         when "00110110101" => index <= 5;
         when "00110110110" => index <= 6;
         when "00110110111" => index <= 5;
         when "00110111000" => index <= 6;
         when "00110111001" => index <= 6;
         when "00110111010" => index <= 6;
         when "00110111011" => index <= 5;
         when "00110111100" => index <= 6;
         when "00110111101" => index <= 5;
         when "00110111110" => index <= 5;
         when "00110111111" => index <= 5;
         when "00111000000" => index <= 8;
         when "00111000001" => index <= 6;
         when "00111000010" => index <= 6;
         when "00111000011" => index <= 5;
         when "00111000100" => index <= 7;
         when "00111000101" => index <= 6;
         when "00111000110" => index <= 6;
         when "00111000111" => index <= 5;
         when "00111001000" => index <= 7;
         when "00111001001" => index <= 6;
         when "00111001010" => index <= 6;
         when "00111001011" => index <= 5;
         when "00111001100" => index <= 6;
         when "00111001101" => index <= 5;
         when "00111001110" => index <= 6;
         when "00111001111" => index <= 5;
         when "00111010000" => index <= 7;
         when "00111010001" => index <= 6;
         when "00111010010" => index <= 6;
         when "00111010011" => index <= 5;
         when "00111010100" => index <= 6;
         when "00111010101" => index <= 6;
         when "00111010110" => index <= 6;
         when "00111010111" => index <= 5;
         when "00111011000" => index <= 7;
         when "00111011001" => index <= 6;
         when "00111011010" => index <= 6;
         when "00111011011" => index <= 5;
         when "00111011100" => index <= 6;
         when "00111011101" => index <= 5;
         when "00111011110" => index <= 5;
         when "00111011111" => index <= 5;
         when "00111100000" => index <= 8;
         when "00111100001" => index <= 6;
         when "00111100010" => index <= 6;
         when "00111100011" => index <= 6;
         when "00111100100" => index <= 7;
         when "00111100101" => index <= 6;
         when "00111100110" => index <= 6;
         when "00111100111" => index <= 5;
         when "00111101000" => index <= 7;
         when "00111101001" => index <= 6;
         when "00111101010" => index <= 6;
         when "00111101011" => index <= 5;
         when "00111101100" => index <= 6;
         when "00111101101" => index <= 5;
         when "00111101110" => index <= 6;
         when "00111101111" => index <= 5;
         when "00111110000" => index <= 7;
         when "00111110001" => index <= 6;
         when "00111110010" => index <= 6;
         when "00111110011" => index <= 5;
         when "00111110100" => index <= 6;
         when "00111110101" => index <= 6;
         when "00111110110" => index <= 6;
         when "00111110111" => index <= 5;
         when "00111111000" => index <= 6;
         when "00111111001" => index <= 6;
         when "00111111010" => index <= 6;
         when "00111111011" => index <= 5;
         when "00111111100" => index <= 6;
         when "00111111101" => index <= 5;
         when "00111111110" => index <= 6;
         when "00111111111" => index <= 5;
         when "01000000000" => index <= 10;
         when "01000000001" => index <= 6;
         when "01000000010" => index <= 6;
         when "01000000011" => index <= 4;
         when "01000000100" => index <= 6;
         when "01000000101" => index <= 5;
         when "01000000110" => index <= 5;
         when "01000000111" => index <= 4;
         when "01000001000" => index <= 7;
         when "01000001001" => index <= 5;
         when "01000001010" => index <= 5;
         when "01000001011" => index <= 4;
         when "01000001100" => index <= 6;
         when "01000001101" => index <= 4;
         when "01000001110" => index <= 5;
         when "01000001111" => index <= 4;
         when "01000010000" => index <= 8;
         when "01000010001" => index <= 5;
         when "01000010010" => index <= 6;
         when "01000010011" => index <= 4;
         when "01000010100" => index <= 6;
         when "01000010101" => index <= 5;
         when "01000010110" => index <= 5;
         when "01000010111" => index <= 4;
         when "01000011000" => index <= 6;
         when "01000011001" => index <= 5;
         when "01000011010" => index <= 5;
         when "01000011011" => index <= 4;
         when "01000011100" => index <= 6;
         when "01000011101" => index <= 5;
         when "01000011110" => index <= 5;
         when "01000011111" => index <= 4;
         when "01000100000" => index <= 8;
         when "01000100001" => index <= 6;
         when "01000100010" => index <= 6;
         when "01000100011" => index <= 5;
         when "01000100100" => index <= 6;
         when "01000100101" => index <= 5;
         when "01000100110" => index <= 5;
         when "01000100111" => index <= 4;
         when "01000101000" => index <= 7;
         when "01000101001" => index <= 5;
         when "01000101010" => index <= 6;
         when "01000101011" => index <= 5;
         when "01000101100" => index <= 6;
         when "01000101101" => index <= 5;
         when "01000101110" => index <= 5;
         when "01000101111" => index <= 4;
         when "01000110000" => index <= 7;
         when "01000110001" => index <= 6;
         when "01000110010" => index <= 6;
         when "01000110011" => index <= 5;
         when "01000110100" => index <= 6;
         when "01000110101" => index <= 5;
         when "01000110110" => index <= 5;
         when "01000110111" => index <= 4;
         when "01000111000" => index <= 6;
         when "01000111001" => index <= 5;
         when "01000111010" => index <= 5;
         when "01000111011" => index <= 5;
         when "01000111100" => index <= 6;
         when "01000111101" => index <= 5;
         when "01000111110" => index <= 5;
         when "01000111111" => index <= 4;
         when "01001000000" => index <= 8;
         when "01001000001" => index <= 6;
         when "01001000010" => index <= 6;
         when "01001000011" => index <= 5;
         when "01001000100" => index <= 7;
         when "01001000101" => index <= 5;
         when "01001000110" => index <= 6;
         when "01001000111" => index <= 5;
         when "01001001000" => index <= 7;
         when "01001001001" => index <= 6;
         when "01001001010" => index <= 6;
         when "01001001011" => index <= 5;
         when "01001001100" => index <= 6;
         when "01001001101" => index <= 5;
         when "01001001110" => index <= 5;
         when "01001001111" => index <= 4;
         when "01001010000" => index <= 7;
         when "01001010001" => index <= 6;
         when "01001010010" => index <= 6;
         when "01001010011" => index <= 5;
         when "01001010100" => index <= 6;
         when "01001010101" => index <= 5;
         when "01001010110" => index <= 5;
         when "01001010111" => index <= 5;
         when "01001011000" => index <= 6;
         when "01001011001" => index <= 5;
         when "01001011010" => index <= 6;
         when "01001011011" => index <= 5;
         when "01001011100" => index <= 6;
         when "01001011101" => index <= 5;
         when "01001011110" => index <= 5;
         when "01001011111" => index <= 5;
         when "01001100000" => index <= 8;
         when "01001100001" => index <= 6;
         when "01001100010" => index <= 6;
         when "01001100011" => index <= 5;
         when "01001100100" => index <= 6;
         when "01001100101" => index <= 5;
         when "01001100110" => index <= 6;
         when "01001100111" => index <= 5;
         when "01001101000" => index <= 7;
         when "01001101001" => index <= 6;
         when "01001101010" => index <= 6;
         when "01001101011" => index <= 5;
         when "01001101100" => index <= 6;
         when "01001101101" => index <= 5;
         when "01001101110" => index <= 5;
         when "01001101111" => index <= 5;
         when "01001110000" => index <= 7;
         when "01001110001" => index <= 6;
         when "01001110010" => index <= 6;
         when "01001110011" => index <= 5;
         when "01001110100" => index <= 6;
         when "01001110101" => index <= 5;
         when "01001110110" => index <= 6;
         when "01001110111" => index <= 5;
         when "01001111000" => index <= 6;
         when "01001111001" => index <= 6;
         when "01001111010" => index <= 6;
         when "01001111011" => index <= 5;
         when "01001111100" => index <= 6;
         when "01001111101" => index <= 5;
         when "01001111110" => index <= 5;
         when "01001111111" => index <= 5;
         when "01010000000" => index <= 9;
         when "01010000001" => index <= 6;
         when "01010000010" => index <= 7;
         when "01010000011" => index <= 5;
         when "01010000100" => index <= 7;
         when "01010000101" => index <= 6;
         when "01010000110" => index <= 6;
         when "01010000111" => index <= 5;
         when "01010001000" => index <= 7;
         when "01010001001" => index <= 6;
         when "01010001010" => index <= 6;
         when "01010001011" => index <= 5;
         when "01010001100" => index <= 6;
         when "01010001101" => index <= 5;
         when "01010001110" => index <= 5;
         when "01010001111" => index <= 5;
         when "01010010000" => index <= 8;
         when "01010010001" => index <= 6;
         when "01010010010" => index <= 6;
         when "01010010011" => index <= 5;
         when "01010010100" => index <= 6;
         when "01010010101" => index <= 5;
         when "01010010110" => index <= 6;
         when "01010010111" => index <= 5;
         when "01010011000" => index <= 7;
         when "01010011001" => index <= 6;
         when "01010011010" => index <= 6;
         when "01010011011" => index <= 5;
         when "01010011100" => index <= 6;
         when "01010011101" => index <= 5;
         when "01010011110" => index <= 5;
         when "01010011111" => index <= 5;
         when "01010100000" => index <= 8;
         when "01010100001" => index <= 6;
         when "01010100010" => index <= 6;
         when "01010100011" => index <= 5;
         when "01010100100" => index <= 7;
         when "01010100101" => index <= 6;
         when "01010100110" => index <= 6;
         when "01010100111" => index <= 5;
         when "01010101000" => index <= 7;
         when "01010101001" => index <= 6;
         when "01010101010" => index <= 6;
         when "01010101011" => index <= 5;
         when "01010101100" => index <= 6;
         when "01010101101" => index <= 5;
         when "01010101110" => index <= 6;
         when "01010101111" => index <= 5;
         when "01010110000" => index <= 7;
         when "01010110001" => index <= 6;
         when "01010110010" => index <= 6;
         when "01010110011" => index <= 5;
         when "01010110100" => index <= 6;
         when "01010110101" => index <= 6;
         when "01010110110" => index <= 6;
         when "01010110111" => index <= 5;
         when "01010111000" => index <= 7;
         when "01010111001" => index <= 6;
         when "01010111010" => index <= 6;
         when "01010111011" => index <= 5;
         when "01010111100" => index <= 6;
         when "01010111101" => index <= 5;
         when "01010111110" => index <= 5;
         when "01010111111" => index <= 5;
         when "01011000000" => index <= 8;
         when "01011000001" => index <= 6;
         when "01011000010" => index <= 7;
         when "01011000011" => index <= 6;
         when "01011000100" => index <= 7;
         when "01011000101" => index <= 6;
         when "01011000110" => index <= 6;
         when "01011000111" => index <= 5;
         when "01011001000" => index <= 7;
         when "01011001001" => index <= 6;
         when "01011001010" => index <= 6;
         when "01011001011" => index <= 5;
         when "01011001100" => index <= 6;
         when "01011001101" => index <= 6;
         when "01011001110" => index <= 6;
         when "01011001111" => index <= 5;
         when "01011010000" => index <= 8;
         when "01011010001" => index <= 6;
         when "01011010010" => index <= 6;
         when "01011010011" => index <= 6;
         when "01011010100" => index <= 7;
         when "01011010101" => index <= 6;
         when "01011010110" => index <= 6;
         when "01011010111" => index <= 5;
         when "01011011000" => index <= 7;
         when "01011011001" => index <= 6;
         when "01011011010" => index <= 6;
         when "01011011011" => index <= 5;
         when "01011011100" => index <= 6;
         when "01011011101" => index <= 5;
         when "01011011110" => index <= 6;
         when "01011011111" => index <= 5;
         when "01011100000" => index <= 8;
         when "01011100001" => index <= 6;
         when "01011100010" => index <= 7;
         when "01011100011" => index <= 6;
         when "01011100100" => index <= 7;
         when "01011100101" => index <= 6;
         when "01011100110" => index <= 6;
         when "01011100111" => index <= 5;
         when "01011101000" => index <= 7;
         when "01011101001" => index <= 6;
         when "01011101010" => index <= 6;
         when "01011101011" => index <= 5;
         when "01011101100" => index <= 6;
         when "01011101101" => index <= 6;
         when "01011101110" => index <= 6;
         when "01011101111" => index <= 5;
         when "01011110000" => index <= 7;
         when "01011110001" => index <= 6;
         when "01011110010" => index <= 6;
         when "01011110011" => index <= 6;
         when "01011110100" => index <= 6;
         when "01011110101" => index <= 6;
         when "01011110110" => index <= 6;
         when "01011110111" => index <= 5;
         when "01011111000" => index <= 7;
         when "01011111001" => index <= 6;
         when "01011111010" => index <= 6;
         when "01011111011" => index <= 5;
         when "01011111100" => index <= 6;
         when "01011111101" => index <= 6;
         when "01011111110" => index <= 6;
         when "01011111111" => index <= 5;
         when "01100000000" => index <= 10;
         when "01100000001" => index <= 7;
         when "01100000010" => index <= 7;
         when "01100000011" => index <= 6;
         when "01100000100" => index <= 7;
         when "01100000101" => index <= 6;
         when "01100000110" => index <= 6;
         when "01100000111" => index <= 5;
         when "01100001000" => index <= 8;
         when "01100001001" => index <= 6;
         when "01100001010" => index <= 6;
         when "01100001011" => index <= 5;
         when "01100001100" => index <= 6;
         when "01100001101" => index <= 5;
         when "01100001110" => index <= 6;
         when "01100001111" => index <= 5;
         when "01100010000" => index <= 8;
         when "01100010001" => index <= 6;
         when "01100010010" => index <= 6;
         when "01100010011" => index <= 5;
         when "01100010100" => index <= 7;
         when "01100010101" => index <= 6;
         when "01100010110" => index <= 6;
         when "01100010111" => index <= 5;
         when "01100011000" => index <= 7;
         when "01100011001" => index <= 6;
         when "01100011010" => index <= 6;
         when "01100011011" => index <= 5;
         when "01100011100" => index <= 6;
         when "01100011101" => index <= 5;
         when "01100011110" => index <= 6;
         when "01100011111" => index <= 5;
         when "01100100000" => index <= 8;
         when "01100100001" => index <= 6;
         when "01100100010" => index <= 7;
         when "01100100011" => index <= 6;
         when "01100100100" => index <= 7;
         when "01100100101" => index <= 6;
         when "01100100110" => index <= 6;
         when "01100100111" => index <= 5;
         when "01100101000" => index <= 7;
         when "01100101001" => index <= 6;
         when "01100101010" => index <= 6;
         when "01100101011" => index <= 5;
         when "01100101100" => index <= 6;
         when "01100101101" => index <= 6;
         when "01100101110" => index <= 6;
         when "01100101111" => index <= 5;
         when "01100110000" => index <= 8;
         when "01100110001" => index <= 6;
         when "01100110010" => index <= 6;
         when "01100110011" => index <= 6;
         when "01100110100" => index <= 7;
         when "01100110101" => index <= 6;
         when "01100110110" => index <= 6;
         when "01100110111" => index <= 5;
         when "01100111000" => index <= 7;
         when "01100111001" => index <= 6;
         when "01100111010" => index <= 6;
         when "01100111011" => index <= 5;
         when "01100111100" => index <= 6;
         when "01100111101" => index <= 5;
         when "01100111110" => index <= 6;
         when "01100111111" => index <= 5;
         when "01101000000" => index <= 9;
         when "01101000001" => index <= 7;
         when "01101000010" => index <= 7;
         when "01101000011" => index <= 6;
         when "01101000100" => index <= 7;
         when "01101000101" => index <= 6;
         when "01101000110" => index <= 6;
         when "01101000111" => index <= 5;
         when "01101001000" => index <= 8;
         when "01101001001" => index <= 6;
         when "01101001010" => index <= 6;
         when "01101001011" => index <= 6;
         when "01101001100" => index <= 7;
         when "01101001101" => index <= 6;
         when "01101001110" => index <= 6;
         when "01101001111" => index <= 5;
         when "01101010000" => index <= 8;
         when "01101010001" => index <= 6;
         when "01101010010" => index <= 7;
         when "01101010011" => index <= 6;
         when "01101010100" => index <= 7;
         when "01101010101" => index <= 6;
         when "01101010110" => index <= 6;
         when "01101010111" => index <= 5;
         when "01101011000" => index <= 7;
         when "01101011001" => index <= 6;
         when "01101011010" => index <= 6;
         when "01101011011" => index <= 5;
         when "01101011100" => index <= 6;
         when "01101011101" => index <= 6;
         when "01101011110" => index <= 6;
         when "01101011111" => index <= 5;
         when "01101100000" => index <= 8;
         when "01101100001" => index <= 7;
         when "01101100010" => index <= 7;
         when "01101100011" => index <= 6;
         when "01101100100" => index <= 7;
         when "01101100101" => index <= 6;
         when "01101100110" => index <= 6;
         when "01101100111" => index <= 5;
         when "01101101000" => index <= 7;
         when "01101101001" => index <= 6;
         when "01101101010" => index <= 6;
         when "01101101011" => index <= 6;
         when "01101101100" => index <= 6;
         when "01101101101" => index <= 6;
         when "01101101110" => index <= 6;
         when "01101101111" => index <= 5;
         when "01101110000" => index <= 7;
         when "01101110001" => index <= 6;
         when "01101110010" => index <= 6;
         when "01101110011" => index <= 6;
         when "01101110100" => index <= 7;
         when "01101110101" => index <= 6;
         when "01101110110" => index <= 6;
         when "01101110111" => index <= 5;
         when "01101111000" => index <= 7;
         when "01101111001" => index <= 6;
         when "01101111010" => index <= 6;
         when "01101111011" => index <= 6;
         when "01101111100" => index <= 6;
         when "01101111101" => index <= 6;
         when "01101111110" => index <= 6;
         when "01101111111" => index <= 5;
         when "01110000000" => index <= 9;
         when "01110000001" => index <= 7;
         when "01110000010" => index <= 7;
         when "01110000011" => index <= 6;
         when "01110000100" => index <= 8;
         when "01110000101" => index <= 6;
         when "01110000110" => index <= 6;
         when "01110000111" => index <= 6;
         when "01110001000" => index <= 8;
         when "01110001001" => index <= 6;
         when "01110001010" => index <= 7;
         when "01110001011" => index <= 6;
         when "01110001100" => index <= 7;
         when "01110001101" => index <= 6;
         when "01110001110" => index <= 6;
         when "01110001111" => index <= 5;
         when "01110010000" => index <= 8;
         when "01110010001" => index <= 7;
         when "01110010010" => index <= 7;
         when "01110010011" => index <= 6;
         when "01110010100" => index <= 7;
         when "01110010101" => index <= 6;
         when "01110010110" => index <= 6;
         when "01110010111" => index <= 5;
         when "01110011000" => index <= 7;
         when "01110011001" => index <= 6;
         when "01110011010" => index <= 6;
         when "01110011011" => index <= 6;
         when "01110011100" => index <= 6;
         when "01110011101" => index <= 6;
         when "01110011110" => index <= 6;
         when "01110011111" => index <= 5;
         when "01110100000" => index <= 8;
         when "01110100001" => index <= 7;
         when "01110100010" => index <= 7;
         when "01110100011" => index <= 6;
         when "01110100100" => index <= 7;
         when "01110100101" => index <= 6;
         when "01110100110" => index <= 6;
         when "01110100111" => index <= 6;
         when "01110101000" => index <= 7;
         when "01110101001" => index <= 6;
         when "01110101010" => index <= 6;
         when "01110101011" => index <= 6;
         when "01110101100" => index <= 7;
         when "01110101101" => index <= 6;
         when "01110101110" => index <= 6;
         when "01110101111" => index <= 5;
         when "01110110000" => index <= 8;
         when "01110110001" => index <= 6;
         when "01110110010" => index <= 7;
         when "01110110011" => index <= 6;
         when "01110110100" => index <= 7;
         when "01110110101" => index <= 6;
         when "01110110110" => index <= 6;
         when "01110110111" => index <= 6;
         when "01110111000" => index <= 7;
         when "01110111001" => index <= 6;
         when "01110111010" => index <= 6;
         when "01110111011" => index <= 6;
         when "01110111100" => index <= 6;
         when "01110111101" => index <= 6;
         when "01110111110" => index <= 6;
         when "01110111111" => index <= 5;
         when "01111000000" => index <= 8;
         when "01111000001" => index <= 7;
         when "01111000010" => index <= 7;
         when "01111000011" => index <= 6;
         when "01111000100" => index <= 7;
         when "01111000101" => index <= 6;
         when "01111000110" => index <= 6;
         when "01111000111" => index <= 6;
         when "01111001000" => index <= 8;
         when "01111001001" => index <= 6;
         when "01111001010" => index <= 7;
         when "01111001011" => index <= 6;
         when "01111001100" => index <= 7;
         when "01111001101" => index <= 6;
         when "01111001110" => index <= 6;
         when "01111001111" => index <= 6;
         when "01111010000" => index <= 8;
         when "01111010001" => index <= 7;
         when "01111010010" => index <= 7;
         when "01111010011" => index <= 6;
         when "01111010100" => index <= 7;
         when "01111010101" => index <= 6;
         when "01111010110" => index <= 6;
         when "01111010111" => index <= 6;
         when "01111011000" => index <= 7;
         when "01111011001" => index <= 6;
         when "01111011010" => index <= 6;
         when "01111011011" => index <= 6;
         when "01111011100" => index <= 7;
         when "01111011101" => index <= 6;
         when "01111011110" => index <= 6;
         when "01111011111" => index <= 5;
         when "01111100000" => index <= 8;
         when "01111100001" => index <= 7;
         when "01111100010" => index <= 7;
         when "01111100011" => index <= 6;
         when "01111100100" => index <= 7;
         when "01111100101" => index <= 6;
         when "01111100110" => index <= 6;
         when "01111100111" => index <= 6;
         when "01111101000" => index <= 7;
         when "01111101001" => index <= 6;
         when "01111101010" => index <= 7;
         when "01111101011" => index <= 6;
         when "01111101100" => index <= 7;
         when "01111101101" => index <= 6;
         when "01111101110" => index <= 6;
         when "01111101111" => index <= 6;
         when "01111110000" => index <= 8;
         when "01111110001" => index <= 7;
         when "01111110010" => index <= 7;
         when "01111110011" => index <= 6;
         when "01111110100" => index <= 7;
         when "01111110101" => index <= 6;
         when "01111110110" => index <= 6;
         when "01111110111" => index <= 6;
         when "01111111000" => index <= 7;
         when "01111111001" => index <= 6;
         when "01111111010" => index <= 6;
         when "01111111011" => index <= 6;
         when "01111111100" => index <= 6;
         when "01111111101" => index <= 6;
         when "01111111110" => index <= 6;
         when "01111111111" => index <= 6;
         when "10000000000" => index <= 11;
         when "10000000001" => index <= 6;
         when "10000000010" => index <= 6;
         when "10000000011" => index <= 5;
         when "10000000100" => index <= 7;
         when "10000000101" => index <= 5;
         when "10000000110" => index <= 5;
         when "10000000111" => index <= 4;
         when "10000001000" => index <= 8;
         when "10000001001" => index <= 5;
         when "10000001010" => index <= 6;
         when "10000001011" => index <= 4;
         when "10000001100" => index <= 6;
         when "10000001101" => index <= 5;
         when "10000001110" => index <= 5;
         when "10000001111" => index <= 4;
         when "10000010000" => index <= 8;
         when "10000010001" => index <= 6;
         when "10000010010" => index <= 6;
         when "10000010011" => index <= 5;
         when "10000010100" => index <= 6;
         when "10000010101" => index <= 5;
         when "10000010110" => index <= 5;
         when "10000010111" => index <= 4;
         when "10000011000" => index <= 7;
         when "10000011001" => index <= 5;
         when "10000011010" => index <= 6;
         when "10000011011" => index <= 5;
         when "10000011100" => index <= 6;
         when "10000011101" => index <= 5;
         when "10000011110" => index <= 5;
         when "10000011111" => index <= 4;
         when "10000100000" => index <= 8;
         when "10000100001" => index <= 6;
         when "10000100010" => index <= 6;
         when "10000100011" => index <= 5;
         when "10000100100" => index <= 7;
         when "10000100101" => index <= 5;
         when "10000100110" => index <= 6;
         when "10000100111" => index <= 5;
         when "10000101000" => index <= 7;
         when "10000101001" => index <= 6;
         when "10000101010" => index <= 6;
         when "10000101011" => index <= 5;
         when "10000101100" => index <= 6;
         when "10000101101" => index <= 5;
         when "10000101110" => index <= 5;
         when "10000101111" => index <= 4;
         when "10000110000" => index <= 7;
         when "10000110001" => index <= 6;
         when "10000110010" => index <= 6;
         when "10000110011" => index <= 5;
         when "10000110100" => index <= 6;
         when "10000110101" => index <= 5;
         when "10000110110" => index <= 5;
         when "10000110111" => index <= 5;
         when "10000111000" => index <= 6;
         when "10000111001" => index <= 5;
         when "10000111010" => index <= 6;
         when "10000111011" => index <= 5;
         when "10000111100" => index <= 6;
         when "10000111101" => index <= 5;
         when "10000111110" => index <= 5;
         when "10000111111" => index <= 5;
         when "10001000000" => index <= 9;
         when "10001000001" => index <= 6;
         when "10001000010" => index <= 7;
         when "10001000011" => index <= 5;
         when "10001000100" => index <= 7;
         when "10001000101" => index <= 6;
         when "10001000110" => index <= 6;
         when "10001000111" => index <= 5;
         when "10001001000" => index <= 7;
         when "10001001001" => index <= 6;
         when "10001001010" => index <= 6;
         when "10001001011" => index <= 5;
         when "10001001100" => index <= 6;
         when "10001001101" => index <= 5;
         when "10001001110" => index <= 5;
         when "10001001111" => index <= 5;
         when "10001010000" => index <= 8;
         when "10001010001" => index <= 6;
         when "10001010010" => index <= 6;
         when "10001010011" => index <= 5;
         when "10001010100" => index <= 6;
         when "10001010101" => index <= 5;
         when "10001010110" => index <= 6;
         when "10001010111" => index <= 5;
         when "10001011000" => index <= 7;
         when "10001011001" => index <= 6;
         when "10001011010" => index <= 6;
         when "10001011011" => index <= 5;
         when "10001011100" => index <= 6;
         when "10001011101" => index <= 5;
         when "10001011110" => index <= 5;
         when "10001011111" => index <= 5;
         when "10001100000" => index <= 8;
         when "10001100001" => index <= 6;
         when "10001100010" => index <= 6;
         when "10001100011" => index <= 5;
         when "10001100100" => index <= 7;
         when "10001100101" => index <= 6;
         when "10001100110" => index <= 6;
         when "10001100111" => index <= 5;
         when "10001101000" => index <= 7;
         when "10001101001" => index <= 6;
         when "10001101010" => index <= 6;
         when "10001101011" => index <= 5;
         when "10001101100" => index <= 6;
         when "10001101101" => index <= 5;
         when "10001101110" => index <= 6;
         when "10001101111" => index <= 5;
         when "10001110000" => index <= 7;
         when "10001110001" => index <= 6;
         when "10001110010" => index <= 6;
         when "10001110011" => index <= 5;
         when "10001110100" => index <= 6;
         when "10001110101" => index <= 6;
         when "10001110110" => index <= 6;
         when "10001110111" => index <= 5;
         when "10001111000" => index <= 7;
         when "10001111001" => index <= 6;
         when "10001111010" => index <= 6;
         when "10001111011" => index <= 5;
         when "10001111100" => index <= 6;
         when "10001111101" => index <= 5;
         when "10001111110" => index <= 5;
         when "10001111111" => index <= 5;
         when "10010000000" => index <= 10;
         when "10010000001" => index <= 7;
         when "10010000010" => index <= 7;
         when "10010000011" => index <= 6;
         when "10010000100" => index <= 7;
         when "10010000101" => index <= 6;
         when "10010000110" => index <= 6;
         when "10010000111" => index <= 5;
         when "10010001000" => index <= 8;
         when "10010001001" => index <= 6;
         when "10010001010" => index <= 6;
         when "10010001011" => index <= 5;
         when "10010001100" => index <= 6;
         when "10010001101" => index <= 5;
         when "10010001110" => index <= 6;
         when "10010001111" => index <= 5;
         when "10010010000" => index <= 8;
         when "10010010001" => index <= 6;
         when "10010010010" => index <= 6;
         when "10010010011" => index <= 5;
         when "10010010100" => index <= 7;
         when "10010010101" => index <= 6;
         when "10010010110" => index <= 6;
         when "10010010111" => index <= 5;
         when "10010011000" => index <= 7;
         when "10010011001" => index <= 6;
         when "10010011010" => index <= 6;
         when "10010011011" => index <= 5;
         when "10010011100" => index <= 6;
         when "10010011101" => index <= 5;
         when "10010011110" => index <= 6;
         when "10010011111" => index <= 5;
         when "10010100000" => index <= 8;
         when "10010100001" => index <= 6;
         when "10010100010" => index <= 7;
         when "10010100011" => index <= 6;
         when "10010100100" => index <= 7;
         when "10010100101" => index <= 6;
         when "10010100110" => index <= 6;
         when "10010100111" => index <= 5;
         when "10010101000" => index <= 7;
         when "10010101001" => index <= 6;
         when "10010101010" => index <= 6;
         when "10010101011" => index <= 5;
         when "10010101100" => index <= 6;
         when "10010101101" => index <= 6;
         when "10010101110" => index <= 6;
         when "10010101111" => index <= 5;
         when "10010110000" => index <= 8;
         when "10010110001" => index <= 6;
         when "10010110010" => index <= 6;
         when "10010110011" => index <= 6;
         when "10010110100" => index <= 7;
         when "10010110101" => index <= 6;
         when "10010110110" => index <= 6;
         when "10010110111" => index <= 5;
         when "10010111000" => index <= 7;
         when "10010111001" => index <= 6;
         when "10010111010" => index <= 6;
         when "10010111011" => index <= 5;
         when "10010111100" => index <= 6;
         when "10010111101" => index <= 5;
         when "10010111110" => index <= 6;
         when "10010111111" => index <= 5;
         when "10011000000" => index <= 9;
         when "10011000001" => index <= 7;
         when "10011000010" => index <= 7;
         when "10011000011" => index <= 6;
         when "10011000100" => index <= 7;
         when "10011000101" => index <= 6;
         when "10011000110" => index <= 6;
         when "10011000111" => index <= 5;
         when "10011001000" => index <= 8;
         when "10011001001" => index <= 6;
         when "10011001010" => index <= 6;
         when "10011001011" => index <= 6;
         when "10011001100" => index <= 7;
         when "10011001101" => index <= 6;
         when "10011001110" => index <= 6;
         when "10011001111" => index <= 5;
         when "10011010000" => index <= 8;
         when "10011010001" => index <= 6;
         when "10011010010" => index <= 7;
         when "10011010011" => index <= 6;
         when "10011010100" => index <= 7;
         when "10011010101" => index <= 6;
         when "10011010110" => index <= 6;
         when "10011010111" => index <= 5;
         when "10011011000" => index <= 7;
         when "10011011001" => index <= 6;
         when "10011011010" => index <= 6;
         when "10011011011" => index <= 5;
         when "10011011100" => index <= 6;
         when "10011011101" => index <= 6;
         when "10011011110" => index <= 6;
         when "10011011111" => index <= 5;
         when "10011100000" => index <= 8;
         when "10011100001" => index <= 7;
         when "10011100010" => index <= 7;
         when "10011100011" => index <= 6;
         when "10011100100" => index <= 7;
         when "10011100101" => index <= 6;
         when "10011100110" => index <= 6;
         when "10011100111" => index <= 5;
         when "10011101000" => index <= 7;
         when "10011101001" => index <= 6;
         when "10011101010" => index <= 6;
         when "10011101011" => index <= 6;
         when "10011101100" => index <= 6;
         when "10011101101" => index <= 6;
         when "10011101110" => index <= 6;
         when "10011101111" => index <= 5;
         when "10011110000" => index <= 7;
         when "10011110001" => index <= 6;
         when "10011110010" => index <= 6;
         when "10011110011" => index <= 6;
         when "10011110100" => index <= 7;
         when "10011110101" => index <= 6;
         when "10011110110" => index <= 6;
         when "10011110111" => index <= 5;
         when "10011111000" => index <= 7;
         when "10011111001" => index <= 6;
         when "10011111010" => index <= 6;
         when "10011111011" => index <= 6;
         when "10011111100" => index <= 6;
         when "10011111101" => index <= 6;
         when "10011111110" => index <= 6;
         when "10011111111" => index <= 5;
         when "10100000000" => index <= 10;
         when "10100000001" => index <= 7;
         when "10100000010" => index <= 7;
         when "10100000011" => index <= 6;
         when "10100000100" => index <= 8;
         when "10100000101" => index <= 6;
         when "10100000110" => index <= 6;
         when "10100000111" => index <= 5;
         when "10100001000" => index <= 8;
         when "10100001001" => index <= 6;
         when "10100001010" => index <= 6;
         when "10100001011" => index <= 5;
         when "10100001100" => index <= 7;
         when "10100001101" => index <= 6;
         when "10100001110" => index <= 6;
         when "10100001111" => index <= 5;
         when "10100010000" => index <= 8;
         when "10100010001" => index <= 6;
         when "10100010010" => index <= 7;
         when "10100010011" => index <= 6;
         when "10100010100" => index <= 7;
         when "10100010101" => index <= 6;
         when "10100010110" => index <= 6;
         when "10100010111" => index <= 5;
         when "10100011000" => index <= 7;
         when "10100011001" => index <= 6;
         when "10100011010" => index <= 6;
         when "10100011011" => index <= 5;
         when "10100011100" => index <= 6;
         when "10100011101" => index <= 6;
         when "10100011110" => index <= 6;
         when "10100011111" => index <= 5;
         when "10100100000" => index <= 9;
         when "10100100001" => index <= 7;
         when "10100100010" => index <= 7;
         when "10100100011" => index <= 6;
         when "10100100100" => index <= 7;
         when "10100100101" => index <= 6;
         when "10100100110" => index <= 6;
         when "10100100111" => index <= 5;
         when "10100101000" => index <= 8;
         when "10100101001" => index <= 6;
         when "10100101010" => index <= 6;
         when "10100101011" => index <= 6;
         when "10100101100" => index <= 7;
         when "10100101101" => index <= 6;
         when "10100101110" => index <= 6;
         when "10100101111" => index <= 5;
         when "10100110000" => index <= 8;
         when "10100110001" => index <= 6;
         when "10100110010" => index <= 7;
         when "10100110011" => index <= 6;
         when "10100110100" => index <= 7;
         when "10100110101" => index <= 6;
         when "10100110110" => index <= 6;
         when "10100110111" => index <= 5;
         when "10100111000" => index <= 7;
         when "10100111001" => index <= 6;
         when "10100111010" => index <= 6;
         when "10100111011" => index <= 5;
         when "10100111100" => index <= 6;
         when "10100111101" => index <= 6;
         when "10100111110" => index <= 6;
         when "10100111111" => index <= 5;
         when "10101000000" => index <= 9;
         when "10101000001" => index <= 7;
         when "10101000010" => index <= 7;
         when "10101000011" => index <= 6;
         when "10101000100" => index <= 8;
         when "10101000101" => index <= 6;
         when "10101000110" => index <= 6;
         when "10101000111" => index <= 6;
         when "10101001000" => index <= 8;
         when "10101001001" => index <= 6;
         when "10101001010" => index <= 7;
         when "10101001011" => index <= 6;
         when "10101001100" => index <= 7;
         when "10101001101" => index <= 6;
         when "10101001110" => index <= 6;
         when "10101001111" => index <= 5;
         when "10101010000" => index <= 8;
         when "10101010001" => index <= 7;
         when "10101010010" => index <= 7;
         when "10101010011" => index <= 6;
         when "10101010100" => index <= 7;
         when "10101010101" => index <= 6;
         when "10101010110" => index <= 6;
         when "10101010111" => index <= 5;
         when "10101011000" => index <= 7;
         when "10101011001" => index <= 6;
         when "10101011010" => index <= 6;
         when "10101011011" => index <= 6;
         when "10101011100" => index <= 6;
         when "10101011101" => index <= 6;
         when "10101011110" => index <= 6;
         when "10101011111" => index <= 5;
         when "10101100000" => index <= 8;
         when "10101100001" => index <= 7;
         when "10101100010" => index <= 7;
         when "10101100011" => index <= 6;
         when "10101100100" => index <= 7;
         when "10101100101" => index <= 6;
         when "10101100110" => index <= 6;
         when "10101100111" => index <= 6;
         when "10101101000" => index <= 7;
         when "10101101001" => index <= 6;
         when "10101101010" => index <= 6;
         when "10101101011" => index <= 6;
         when "10101101100" => index <= 7;
         when "10101101101" => index <= 6;
         when "10101101110" => index <= 6;
         when "10101101111" => index <= 5;
         when "10101110000" => index <= 8;
         when "10101110001" => index <= 6;
         when "10101110010" => index <= 7;
         when "10101110011" => index <= 6;
         when "10101110100" => index <= 7;
         when "10101110101" => index <= 6;
         when "10101110110" => index <= 6;
         when "10101110111" => index <= 6;
         when "10101111000" => index <= 7;
         when "10101111001" => index <= 6;
         when "10101111010" => index <= 6;
         when "10101111011" => index <= 6;
         when "10101111100" => index <= 6;
         when "10101111101" => index <= 6;
         when "10101111110" => index <= 6;
         when "10101111111" => index <= 5;
         when "10110000000" => index <= 9;
         when "10110000001" => index <= 7;
         when "10110000010" => index <= 8;
         when "10110000011" => index <= 6;
         when "10110000100" => index <= 8;
         when "10110000101" => index <= 6;
         when "10110000110" => index <= 7;
         when "10110000111" => index <= 6;
         when "10110001000" => index <= 8;
         when "10110001001" => index <= 7;
         when "10110001010" => index <= 7;
         when "10110001011" => index <= 6;
         when "10110001100" => index <= 7;
         when "10110001101" => index <= 6;
         when "10110001110" => index <= 6;
         when "10110001111" => index <= 5;
         when "10110010000" => index <= 8;
         when "10110010001" => index <= 7;
         when "10110010010" => index <= 7;
         when "10110010011" => index <= 6;
         when "10110010100" => index <= 7;
         when "10110010101" => index <= 6;
         when "10110010110" => index <= 6;
         when "10110010111" => index <= 6;
         when "10110011000" => index <= 7;
         when "10110011001" => index <= 6;
         when "10110011010" => index <= 6;
         when "10110011011" => index <= 6;
         when "10110011100" => index <= 7;
         when "10110011101" => index <= 6;
         when "10110011110" => index <= 6;
         when "10110011111" => index <= 5;
         when "10110100000" => index <= 8;
         when "10110100001" => index <= 7;
         when "10110100010" => index <= 7;
         when "10110100011" => index <= 6;
         when "10110100100" => index <= 7;
         when "10110100101" => index <= 6;
         when "10110100110" => index <= 6;
         when "10110100111" => index <= 6;
         when "10110101000" => index <= 8;
         when "10110101001" => index <= 6;
         when "10110101010" => index <= 7;
         when "10110101011" => index <= 6;
         when "10110101100" => index <= 7;
         when "10110101101" => index <= 6;
         when "10110101110" => index <= 6;
         when "10110101111" => index <= 6;
         when "10110110000" => index <= 8;
         when "10110110001" => index <= 7;
         when "10110110010" => index <= 7;
         when "10110110011" => index <= 6;
         when "10110110100" => index <= 7;
         when "10110110101" => index <= 6;
         when "10110110110" => index <= 6;
         when "10110110111" => index <= 6;
         when "10110111000" => index <= 7;
         when "10110111001" => index <= 6;
         when "10110111010" => index <= 6;
         when "10110111011" => index <= 6;
         when "10110111100" => index <= 7;
         when "10110111101" => index <= 6;
         when "10110111110" => index <= 6;
         when "10110111111" => index <= 5;
         when "10111000000" => index <= 9;
         when "10111000001" => index <= 7;
         when "10111000010" => index <= 7;
         when "10111000011" => index <= 6;
         when "10111000100" => index <= 8;
         when "10111000101" => index <= 6;
         when "10111000110" => index <= 7;
         when "10111000111" => index <= 6;
         when "10111001000" => index <= 8;
         when "10111001001" => index <= 7;
         when "10111001010" => index <= 7;
         when "10111001011" => index <= 6;
         when "10111001100" => index <= 7;
         when "10111001101" => index <= 6;
         when "10111001110" => index <= 6;
         when "10111001111" => index <= 6;
         when "10111010000" => index <= 8;
         when "10111010001" => index <= 7;
         when "10111010010" => index <= 7;
         when "10111010011" => index <= 6;
         when "10111010100" => index <= 7;
         when "10111010101" => index <= 6;
         when "10111010110" => index <= 6;
         when "10111010111" => index <= 6;
         when "10111011000" => index <= 7;
         when "10111011001" => index <= 6;
         when "10111011010" => index <= 7;
         when "10111011011" => index <= 6;
         when "10111011100" => index <= 7;
         when "10111011101" => index <= 6;
         when "10111011110" => index <= 6;
         when "10111011111" => index <= 6;
         when "10111100000" => index <= 8;
         when "10111100001" => index <= 7;
         when "10111100010" => index <= 7;
         when "10111100011" => index <= 6;
         when "10111100100" => index <= 7;
         when "10111100101" => index <= 6;
         when "10111100110" => index <= 7;
         when "10111100111" => index <= 6;
         when "10111101000" => index <= 8;
         when "10111101001" => index <= 7;
         when "10111101010" => index <= 7;
         when "10111101011" => index <= 6;
         when "10111101100" => index <= 7;
         when "10111101101" => index <= 6;
         when "10111101110" => index <= 6;
         when "10111101111" => index <= 6;
         when "10111110000" => index <= 8;
         when "10111110001" => index <= 7;
         when "10111110010" => index <= 7;
         when "10111110011" => index <= 6;
         when "10111110100" => index <= 7;
         when "10111110101" => index <= 6;
         when "10111110110" => index <= 6;
         when "10111110111" => index <= 6;
         when "10111111000" => index <= 7;
         when "10111111001" => index <= 6;
         when "10111111010" => index <= 6;
         when "10111111011" => index <= 6;
         when "10111111100" => index <= 7;
         when "10111111101" => index <= 6;
         when "10111111110" => index <= 6;
         when "10111111111" => index <= 6;
         when "11000000000" => index <= 10;
         when "11000000001" => index <= 7;
         when "11000000010" => index <= 8;
         when "11000000011" => index <= 6;
         when "11000000100" => index <= 8;
         when "11000000101" => index <= 6;
         when "11000000110" => index <= 6;
         when "11000000111" => index <= 5;
         when "11000001000" => index <= 8;
         when "11000001001" => index <= 6;
         when "11000001010" => index <= 7;
         when "11000001011" => index <= 6;
         when "11000001100" => index <= 7;
         when "11000001101" => index <= 6;
         when "11000001110" => index <= 6;
         when "11000001111" => index <= 5;
         when "11000010000" => index <= 9;
         when "11000010001" => index <= 7;
         when "11000010010" => index <= 7;
         when "11000010011" => index <= 6;
         when "11000010100" => index <= 7;
         when "11000010101" => index <= 6;
         when "11000010110" => index <= 6;
         when "11000010111" => index <= 5;
         when "11000011000" => index <= 8;
         when "11000011001" => index <= 6;
         when "11000011010" => index <= 6;
         when "11000011011" => index <= 6;
         when "11000011100" => index <= 7;
         when "11000011101" => index <= 6;
         when "11000011110" => index <= 6;
         when "11000011111" => index <= 5;
         when "11000100000" => index <= 9;
         when "11000100001" => index <= 7;
         when "11000100010" => index <= 7;
         when "11000100011" => index <= 6;
         when "11000100100" => index <= 8;
         when "11000100101" => index <= 6;
         when "11000100110" => index <= 6;
         when "11000100111" => index <= 6;
         when "11000101000" => index <= 8;
         when "11000101001" => index <= 6;
         when "11000101010" => index <= 7;
         when "11000101011" => index <= 6;
         when "11000101100" => index <= 7;
         when "11000101101" => index <= 6;
         when "11000101110" => index <= 6;
         when "11000101111" => index <= 5;
         when "11000110000" => index <= 8;
         when "11000110001" => index <= 7;
         when "11000110010" => index <= 7;
         when "11000110011" => index <= 6;
         when "11000110100" => index <= 7;
         when "11000110101" => index <= 6;
         when "11000110110" => index <= 6;
         when "11000110111" => index <= 5;
         when "11000111000" => index <= 7;
         when "11000111001" => index <= 6;
         when "11000111010" => index <= 6;
         when "11000111011" => index <= 6;
         when "11000111100" => index <= 6;
         when "11000111101" => index <= 6;
         when "11000111110" => index <= 6;
         when "11000111111" => index <= 5;
         when "11001000000" => index <= 9;
         when "11001000001" => index <= 7;
         when "11001000010" => index <= 8;
         when "11001000011" => index <= 6;
         when "11001000100" => index <= 8;
         when "11001000101" => index <= 6;
         when "11001000110" => index <= 7;
         when "11001000111" => index <= 6;
         when "11001001000" => index <= 8;
         when "11001001001" => index <= 7;
         when "11001001010" => index <= 7;
         when "11001001011" => index <= 6;
         when "11001001100" => index <= 7;
         when "11001001101" => index <= 6;
         when "11001001110" => index <= 6;
         when "11001001111" => index <= 5;
         when "11001010000" => index <= 8;
         when "11001010001" => index <= 7;
         when "11001010010" => index <= 7;
         when "11001010011" => index <= 6;
         when "11001010100" => index <= 7;
         when "11001010101" => index <= 6;
         when "11001010110" => index <= 6;
         when "11001010111" => index <= 6;
         when "11001011000" => index <= 7;
         when "11001011001" => index <= 6;
         when "11001011010" => index <= 6;
         when "11001011011" => index <= 6;
         when "11001011100" => index <= 7;
         when "11001011101" => index <= 6;
         when "11001011110" => index <= 6;
         when "11001011111" => index <= 5;
         when "11001100000" => index <= 8;
         when "11001100001" => index <= 7;
         when "11001100010" => index <= 7;
         when "11001100011" => index <= 6;
         when "11001100100" => index <= 7;
         when "11001100101" => index <= 6;
         when "11001100110" => index <= 6;
         when "11001100111" => index <= 6;
         when "11001101000" => index <= 8;
         when "11001101001" => index <= 6;
         when "11001101010" => index <= 7;
         when "11001101011" => index <= 6;
         when "11001101100" => index <= 7;
         when "11001101101" => index <= 6;
         when "11001101110" => index <= 6;
         when "11001101111" => index <= 6;
         when "11001110000" => index <= 8;
         when "11001110001" => index <= 7;
         when "11001110010" => index <= 7;
         when "11001110011" => index <= 6;
         when "11001110100" => index <= 7;
         when "11001110101" => index <= 6;
         when "11001110110" => index <= 6;
         when "11001110111" => index <= 6;
         when "11001111000" => index <= 7;
         when "11001111001" => index <= 6;
         when "11001111010" => index <= 6;
         when "11001111011" => index <= 6;
         when "11001111100" => index <= 7;
         when "11001111101" => index <= 6;
         when "11001111110" => index <= 6;
         when "11001111111" => index <= 5;
         when "11010000000" => index <= 10;
         when "11010000001" => index <= 8;
         when "11010000010" => index <= 8;
         when "11010000011" => index <= 6;
         when "11010000100" => index <= 8;
         when "11010000101" => index <= 7;
         when "11010000110" => index <= 7;
         when "11010000111" => index <= 6;
         when "11010001000" => index <= 8;
         when "11010001001" => index <= 7;
         when "11010001010" => index <= 7;
         when "11010001011" => index <= 6;
         when "11010001100" => index <= 7;
         when "11010001101" => index <= 6;
         when "11010001110" => index <= 6;
         when "11010001111" => index <= 6;
         when "11010010000" => index <= 8;
         when "11010010001" => index <= 7;
         when "11010010010" => index <= 7;
         when "11010010011" => index <= 6;
         when "11010010100" => index <= 7;
         when "11010010101" => index <= 6;
         when "11010010110" => index <= 6;
         when "11010010111" => index <= 6;
         when "11010011000" => index <= 8;
         when "11010011001" => index <= 6;
         when "11010011010" => index <= 7;
         when "11010011011" => index <= 6;
         when "11010011100" => index <= 7;
         when "11010011101" => index <= 6;
         when "11010011110" => index <= 6;
         when "11010011111" => index <= 6;
         when "11010100000" => index <= 9;
         when "11010100001" => index <= 7;
         when "11010100010" => index <= 7;
         when "11010100011" => index <= 6;
         when "11010100100" => index <= 8;
         when "11010100101" => index <= 6;
         when "11010100110" => index <= 7;
         when "11010100111" => index <= 6;
         when "11010101000" => index <= 8;
         when "11010101001" => index <= 7;
         when "11010101010" => index <= 7;
         when "11010101011" => index <= 6;
         when "11010101100" => index <= 7;
         when "11010101101" => index <= 6;
         when "11010101110" => index <= 6;
         when "11010101111" => index <= 6;
         when "11010110000" => index <= 8;
         when "11010110001" => index <= 7;
         when "11010110010" => index <= 7;
         when "11010110011" => index <= 6;
         when "11010110100" => index <= 7;
         when "11010110101" => index <= 6;
         when "11010110110" => index <= 6;
         when "11010110111" => index <= 6;
         when "11010111000" => index <= 7;
         when "11010111001" => index <= 6;
         when "11010111010" => index <= 7;
         when "11010111011" => index <= 6;
         when "11010111100" => index <= 7;
         when "11010111101" => index <= 6;
         when "11010111110" => index <= 6;
         when "11010111111" => index <= 6;
         when "11011000000" => index <= 9;
         when "11011000001" => index <= 7;
         when "11011000010" => index <= 8;
         when "11011000011" => index <= 6;
         when "11011000100" => index <= 8;
         when "11011000101" => index <= 7;
         when "11011000110" => index <= 7;
         when "11011000111" => index <= 6;
         when "11011001000" => index <= 8;
         when "11011001001" => index <= 7;
         when "11011001010" => index <= 7;
         when "11011001011" => index <= 6;
         when "11011001100" => index <= 7;
         when "11011001101" => index <= 6;
         when "11011001110" => index <= 6;
         when "11011001111" => index <= 6;
         when "11011010000" => index <= 8;
         when "11011010001" => index <= 7;
         when "11011010010" => index <= 7;
         when "11011010011" => index <= 6;
         when "11011010100" => index <= 7;
         when "11011010101" => index <= 6;
         when "11011010110" => index <= 7;
         when "11011010111" => index <= 6;
         when "11011011000" => index <= 8;
         when "11011011001" => index <= 7;
         when "11011011010" => index <= 7;
         when "11011011011" => index <= 6;
         when "11011011100" => index <= 7;
         when "11011011101" => index <= 6;
         when "11011011110" => index <= 6;
         when "11011011111" => index <= 6;
         when "11011100000" => index <= 8;
         when "11011100001" => index <= 7;
         when "11011100010" => index <= 7;
         when "11011100011" => index <= 6;
         when "11011100100" => index <= 8;
         when "11011100101" => index <= 7;
         when "11011100110" => index <= 7;
         when "11011100111" => index <= 6;
         when "11011101000" => index <= 8;
         when "11011101001" => index <= 7;
         when "11011101010" => index <= 7;
         when "11011101011" => index <= 6;
         when "11011101100" => index <= 7;
         when "11011101101" => index <= 6;
         when "11011101110" => index <= 6;
         when "11011101111" => index <= 6;
         when "11011110000" => index <= 8;
         when "11011110001" => index <= 7;
         when "11011110010" => index <= 7;
         when "11011110011" => index <= 6;
         when "11011110100" => index <= 7;
         when "11011110101" => index <= 6;
         when "11011110110" => index <= 6;
         when "11011110111" => index <= 6;
         when "11011111000" => index <= 7;
         when "11011111001" => index <= 6;
         when "11011111010" => index <= 7;
         when "11011111011" => index <= 6;
         when "11011111100" => index <= 7;
         when "11011111101" => index <= 6;
         when "11011111110" => index <= 6;
         when "11011111111" => index <= 6;
         when "11100000000" => index <= 10;
         when "11100000001" => index <= 8;
         when "11100000010" => index <= 8;
         when "11100000011" => index <= 7;
         when "11100000100" => index <= 8;
         when "11100000101" => index <= 7;
         when "11100000110" => index <= 7;
         when "11100000111" => index <= 6;
         when "11100001000" => index <= 8;
         when "11100001001" => index <= 7;
         when "11100001010" => index <= 7;
         when "11100001011" => index <= 6;
         when "11100001100" => index <= 7;
         when "11100001101" => index <= 6;
         when "11100001110" => index <= 6;
         when "11100001111" => index <= 6;
         when "11100010000" => index <= 9;
         when "11100010001" => index <= 7;
         when "11100010010" => index <= 7;
         when "11100010011" => index <= 6;
         when "11100010100" => index <= 8;
         when "11100010101" => index <= 6;
         when "11100010110" => index <= 7;
         when "11100010111" => index <= 6;
         when "11100011000" => index <= 8;
         when "11100011001" => index <= 7;
         when "11100011010" => index <= 7;
         when "11100011011" => index <= 6;
         when "11100011100" => index <= 7;
         when "11100011101" => index <= 6;
         when "11100011110" => index <= 6;
         when "11100011111" => index <= 6;
         when "11100100000" => index <= 9;
         when "11100100001" => index <= 7;
         when "11100100010" => index <= 8;
         when "11100100011" => index <= 6;
         when "11100100100" => index <= 8;
         when "11100100101" => index <= 7;
         when "11100100110" => index <= 7;
         when "11100100111" => index <= 6;
         when "11100101000" => index <= 8;
         when "11100101001" => index <= 7;
         when "11100101010" => index <= 7;
         when "11100101011" => index <= 6;
         when "11100101100" => index <= 7;
         when "11100101101" => index <= 6;
         when "11100101110" => index <= 6;
         when "11100101111" => index <= 6;
         when "11100110000" => index <= 8;
         when "11100110001" => index <= 7;
         when "11100110010" => index <= 7;
         when "11100110011" => index <= 6;
         when "11100110100" => index <= 7;
         when "11100110101" => index <= 6;
         when "11100110110" => index <= 7;
         when "11100110111" => index <= 6;
         when "11100111000" => index <= 8;
         when "11100111001" => index <= 7;
         when "11100111010" => index <= 7;
         when "11100111011" => index <= 6;
         when "11100111100" => index <= 7;
         when "11100111101" => index <= 6;
         when "11100111110" => index <= 6;
         when "11100111111" => index <= 6;
         when "11101000000" => index <= 9;
         when "11101000001" => index <= 8;
         when "11101000010" => index <= 8;
         when "11101000011" => index <= 7;
         when "11101000100" => index <= 8;
         when "11101000101" => index <= 7;
         when "11101000110" => index <= 7;
         when "11101000111" => index <= 6;
         when "11101001000" => index <= 8;
         when "11101001001" => index <= 7;
         when "11101001010" => index <= 7;
         when "11101001011" => index <= 6;
         when "11101001100" => index <= 7;
         when "11101001101" => index <= 6;
         when "11101001110" => index <= 7;
         when "11101001111" => index <= 6;
         when "11101010000" => index <= 8;
         when "11101010001" => index <= 7;
         when "11101010010" => index <= 7;
         when "11101010011" => index <= 6;
         when "11101010100" => index <= 8;
         when "11101010101" => index <= 7;
         when "11101010110" => index <= 7;
         when "11101010111" => index <= 6;
         when "11101011000" => index <= 8;
         when "11101011001" => index <= 7;
         when "11101011010" => index <= 7;
         when "11101011011" => index <= 6;
         when "11101011100" => index <= 7;
         when "11101011101" => index <= 6;
         when "11101011110" => index <= 6;
         when "11101011111" => index <= 6;
         when "11101100000" => index <= 9;
         when "11101100001" => index <= 7;
         when "11101100010" => index <= 8;
         when "11101100011" => index <= 7;
         when "11101100100" => index <= 8;
         when "11101100101" => index <= 7;
         when "11101100110" => index <= 7;
         when "11101100111" => index <= 6;
         when "11101101000" => index <= 8;
         when "11101101001" => index <= 7;
         when "11101101010" => index <= 7;
         when "11101101011" => index <= 6;
         when "11101101100" => index <= 7;
         when "11101101101" => index <= 6;
         when "11101101110" => index <= 6;
         when "11101101111" => index <= 6;
         when "11101110000" => index <= 8;
         when "11101110001" => index <= 7;
         when "11101110010" => index <= 7;
         when "11101110011" => index <= 6;
         when "11101110100" => index <= 7;
         when "11101110101" => index <= 6;
         when "11101110110" => index <= 7;
         when "11101110111" => index <= 6;
         when "11101111000" => index <= 7;
         when "11101111001" => index <= 7;
         when "11101111010" => index <= 7;
         when "11101111011" => index <= 6;
         when "11101111100" => index <= 7;
         when "11101111101" => index <= 6;
         when "11101111110" => index <= 6;
         when "11101111111" => index <= 6;
         when "11110000000" => index <= 10;
         when "11110000001" => index <= 8;
         when "11110000010" => index <= 8;
         when "11110000011" => index <= 7;
         when "11110000100" => index <= 8;
         when "11110000101" => index <= 7;
         when "11110000110" => index <= 7;
         when "11110000111" => index <= 6;
         when "11110001000" => index <= 8;
         when "11110001001" => index <= 7;
         when "11110001010" => index <= 7;
         when "11110001011" => index <= 6;
         when "11110001100" => index <= 8;
         when "11110001101" => index <= 7;
         when "11110001110" => index <= 7;
         when "11110001111" => index <= 6;
         when "11110010000" => index <= 9;
         when "11110010001" => index <= 7;
         when "11110010010" => index <= 8;
         when "11110010011" => index <= 7;
         when "11110010100" => index <= 8;
         when "11110010101" => index <= 7;
         when "11110010110" => index <= 7;
         when "11110010111" => index <= 6;
         when "11110011000" => index <= 8;
         when "11110011001" => index <= 7;
         when "11110011010" => index <= 7;
         when "11110011011" => index <= 6;
         when "11110011100" => index <= 7;
         when "11110011101" => index <= 6;
         when "11110011110" => index <= 6;
         when "11110011111" => index <= 6;
         when "11110100000" => index <= 9;
         when "11110100001" => index <= 8;
         when "11110100010" => index <= 8;
         when "11110100011" => index <= 7;
         when "11110100100" => index <= 8;
         when "11110100101" => index <= 7;
         when "11110100110" => index <= 7;
         when "11110100111" => index <= 6;
         when "11110101000" => index <= 8;
         when "11110101001" => index <= 7;
         when "11110101010" => index <= 7;
         when "11110101011" => index <= 6;
         when "11110101100" => index <= 7;
         when "11110101101" => index <= 6;
         when "11110101110" => index <= 7;
         when "11110101111" => index <= 6;
         when "11110110000" => index <= 8;
         when "11110110001" => index <= 7;
         when "11110110010" => index <= 7;
         when "11110110011" => index <= 6;
         when "11110110100" => index <= 7;
         when "11110110101" => index <= 7;
         when "11110110110" => index <= 7;
         when "11110110111" => index <= 6;
         when "11110111000" => index <= 8;
         when "11110111001" => index <= 7;
         when "11110111010" => index <= 7;
         when "11110111011" => index <= 6;
         when "11110111100" => index <= 7;
         when "11110111101" => index <= 6;
         when "11110111110" => index <= 6;
         when "11110111111" => index <= 6;
         when "11111000000" => index <= 9;
         when "11111000001" => index <= 8;
         when "11111000010" => index <= 8;
         when "11111000011" => index <= 7;
         when "11111000100" => index <= 8;
         when "11111000101" => index <= 7;
         when "11111000110" => index <= 7;
         when "11111000111" => index <= 6;
         when "11111001000" => index <= 8;
         when "11111001001" => index <= 7;
         when "11111001010" => index <= 7;
         when "11111001011" => index <= 6;
         when "11111001100" => index <= 7;
         when "11111001101" => index <= 7;
         when "11111001110" => index <= 7;
         when "11111001111" => index <= 6;
         when "11111010000" => index <= 8;
         when "11111010001" => index <= 7;
         when "11111010010" => index <= 7;
         when "11111010011" => index <= 7;
         when "11111010100" => index <= 8;
         when "11111010101" => index <= 7;
         when "11111010110" => index <= 7;
         when "11111010111" => index <= 6;
         when "11111011000" => index <= 8;
         when "11111011001" => index <= 7;
         when "11111011010" => index <= 7;
         when "11111011011" => index <= 6;
         when "11111011100" => index <= 7;
         when "11111011101" => index <= 6;
         when "11111011110" => index <= 7;
         when "11111011111" => index <= 6;
         when "11111100000" => index <= 8;
         when "11111100001" => index <= 7;
         when "11111100010" => index <= 8;
         when "11111100011" => index <= 7;
         when "11111100100" => index <= 8;
         when "11111100101" => index <= 7;
         when "11111100110" => index <= 7;
         when "11111100111" => index <= 6;
         when "11111101000" => index <= 8;
         when "11111101001" => index <= 7;
         when "11111101010" => index <= 7;
         when "11111101011" => index <= 6;
         when "11111101100" => index <= 7;
         when "11111101101" => index <= 7;
         when "11111101110" => index <= 7;
         when "11111101111" => index <= 6;
         when "11111110000" => index <= 8;
         when "11111110001" => index <= 7;
         when "11111110010" => index <= 7;
         when "11111110011" => index <= 7;
         when "11111110100" => index <= 7;
         when "11111110101" => index <= 7;
         when "11111110110" => index <= 7;
         when "11111110111" => index <= 6;
         when "11111111000" => index <= 8;
         when "11111111001" => index <= 7;
         when "11111111010" => index <= 7;
         when "11111111011" => index <= 6;
         when "11111111100" => index <= 7;
         when "11111111101" => index <= 6;
         when "11111111110" => index <= 6;
         when "11111111111" => index <= 6;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_12 : if (length = 12) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "000000000000" => index <= 0;
         when "000000000001" => index <= 1;
         when "000000000010" => index <= 2;
         when "000000000011" => index <= 2;
         when "000000000100" => index <= 3;
         when "000000000101" => index <= 2;
         when "000000000110" => index <= 2;
         when "000000000111" => index <= 2;
         when "000000001000" => index <= 4;
         when "000000001001" => index <= 2;
         when "000000001010" => index <= 3;
         when "000000001011" => index <= 2;
         when "000000001100" => index <= 4;
         when "000000001101" => index <= 3;
         when "000000001110" => index <= 3;
         when "000000001111" => index <= 2;
         when "000000010000" => index <= 5;
         when "000000010001" => index <= 3;
         when "000000010010" => index <= 4;
         when "000000010011" => index <= 3;
         when "000000010100" => index <= 4;
         when "000000010101" => index <= 3;
         when "000000010110" => index <= 3;
         when "000000010111" => index <= 3;
         when "000000011000" => index <= 4;
         when "000000011001" => index <= 3;
         when "000000011010" => index <= 4;
         when "000000011011" => index <= 3;
         when "000000011100" => index <= 4;
         when "000000011101" => index <= 3;
         when "000000011110" => index <= 4;
         when "000000011111" => index <= 3;
         when "000000100000" => index <= 6;
         when "000000100001" => index <= 4;
         when "000000100010" => index <= 4;
         when "000000100011" => index <= 3;
         when "000000100100" => index <= 4;
         when "000000100101" => index <= 3;
         when "000000100110" => index <= 4;
         when "000000100111" => index <= 3;
         when "000000101000" => index <= 5;
         when "000000101001" => index <= 4;
         when "000000101010" => index <= 4;
         when "000000101011" => index <= 3;
         when "000000101100" => index <= 4;
         when "000000101101" => index <= 4;
         when "000000101110" => index <= 4;
         when "000000101111" => index <= 3;
         when "000000110000" => index <= 6;
         when "000000110001" => index <= 4;
         when "000000110010" => index <= 4;
         when "000000110011" => index <= 4;
         when "000000110100" => index <= 5;
         when "000000110101" => index <= 4;
         when "000000110110" => index <= 4;
         when "000000110111" => index <= 3;
         when "000000111000" => index <= 5;
         when "000000111001" => index <= 4;
         when "000000111010" => index <= 4;
         when "000000111011" => index <= 4;
         when "000000111100" => index <= 4;
         when "000000111101" => index <= 4;
         when "000000111110" => index <= 4;
         when "000000111111" => index <= 4;
         when "000001000000" => index <= 7;
         when "000001000001" => index <= 4;
         when "000001000010" => index <= 4;
         when "000001000011" => index <= 3;
         when "000001000100" => index <= 5;
         when "000001000101" => index <= 4;
         when "000001000110" => index <= 4;
         when "000001000111" => index <= 3;
         when "000001001000" => index <= 6;
         when "000001001001" => index <= 4;
         when "000001001010" => index <= 4;
         when "000001001011" => index <= 4;
         when "000001001100" => index <= 5;
         when "000001001101" => index <= 4;
         when "000001001110" => index <= 4;
         when "000001001111" => index <= 3;
         when "000001010000" => index <= 6;
         when "000001010001" => index <= 4;
         when "000001010010" => index <= 5;
         when "000001010011" => index <= 4;
         when "000001010100" => index <= 5;
         when "000001010101" => index <= 4;
         when "000001010110" => index <= 4;
         when "000001010111" => index <= 4;
         when "000001011000" => index <= 5;
         when "000001011001" => index <= 4;
         when "000001011010" => index <= 4;
         when "000001011011" => index <= 4;
         when "000001011100" => index <= 5;
         when "000001011101" => index <= 4;
         when "000001011110" => index <= 4;
         when "000001011111" => index <= 4;
         when "000001100000" => index <= 6;
         when "000001100001" => index <= 5;
         when "000001100010" => index <= 5;
         when "000001100011" => index <= 4;
         when "000001100100" => index <= 5;
         when "000001100101" => index <= 4;
         when "000001100110" => index <= 4;
         when "000001100111" => index <= 4;
         when "000001101000" => index <= 6;
         when "000001101001" => index <= 4;
         when "000001101010" => index <= 5;
         when "000001101011" => index <= 4;
         when "000001101100" => index <= 5;
         when "000001101101" => index <= 4;
         when "000001101110" => index <= 4;
         when "000001101111" => index <= 4;
         when "000001110000" => index <= 6;
         when "000001110001" => index <= 5;
         when "000001110010" => index <= 5;
         when "000001110011" => index <= 4;
         when "000001110100" => index <= 5;
         when "000001110101" => index <= 4;
         when "000001110110" => index <= 5;
         when "000001110111" => index <= 4;
         when "000001111000" => index <= 6;
         when "000001111001" => index <= 5;
         when "000001111010" => index <= 5;
         when "000001111011" => index <= 4;
         when "000001111100" => index <= 5;
         when "000001111101" => index <= 4;
         when "000001111110" => index <= 4;
         when "000001111111" => index <= 4;
         when "000010000000" => index <= 8;
         when "000010000001" => index <= 4;
         when "000010000010" => index <= 5;
         when "000010000011" => index <= 4;
         when "000010000100" => index <= 6;
         when "000010000101" => index <= 4;
         when "000010000110" => index <= 4;
         when "000010000111" => index <= 4;
         when "000010001000" => index <= 6;
         when "000010001001" => index <= 4;
         when "000010001010" => index <= 5;
         when "000010001011" => index <= 4;
         when "000010001100" => index <= 5;
         when "000010001101" => index <= 4;
         when "000010001110" => index <= 4;
         when "000010001111" => index <= 4;
         when "000010010000" => index <= 6;
         when "000010010001" => index <= 5;
         when "000010010010" => index <= 5;
         when "000010010011" => index <= 4;
         when "000010010100" => index <= 5;
         when "000010010101" => index <= 4;
         when "000010010110" => index <= 4;
         when "000010010111" => index <= 4;
         when "000010011000" => index <= 6;
         when "000010011001" => index <= 4;
         when "000010011010" => index <= 5;
         when "000010011011" => index <= 4;
         when "000010011100" => index <= 5;
         when "000010011101" => index <= 4;
         when "000010011110" => index <= 4;
         when "000010011111" => index <= 4;
         when "000010100000" => index <= 7;
         when "000010100001" => index <= 5;
         when "000010100010" => index <= 5;
         when "000010100011" => index <= 4;
         when "000010100100" => index <= 6;
         when "000010100101" => index <= 4;
         when "000010100110" => index <= 5;
         when "000010100111" => index <= 4;
         when "000010101000" => index <= 6;
         when "000010101001" => index <= 5;
         when "000010101010" => index <= 5;
         when "000010101011" => index <= 4;
         when "000010101100" => index <= 5;
         when "000010101101" => index <= 4;
         when "000010101110" => index <= 5;
         when "000010101111" => index <= 4;
         when "000010110000" => index <= 6;
         when "000010110001" => index <= 5;
         when "000010110010" => index <= 5;
         when "000010110011" => index <= 4;
         when "000010110100" => index <= 6;
         when "000010110101" => index <= 5;
         when "000010110110" => index <= 5;
         when "000010110111" => index <= 4;
         when "000010111000" => index <= 6;
         when "000010111001" => index <= 5;
         when "000010111010" => index <= 5;
         when "000010111011" => index <= 4;
         when "000010111100" => index <= 5;
         when "000010111101" => index <= 4;
         when "000010111110" => index <= 5;
         when "000010111111" => index <= 4;
         when "000011000000" => index <= 8;
         when "000011000001" => index <= 5;
         when "000011000010" => index <= 6;
         when "000011000011" => index <= 4;
         when "000011000100" => index <= 6;
         when "000011000101" => index <= 5;
         when "000011000110" => index <= 5;
         when "000011000111" => index <= 4;
         when "000011001000" => index <= 6;
         when "000011001001" => index <= 5;
         when "000011001010" => index <= 5;
         when "000011001011" => index <= 4;
         when "000011001100" => index <= 6;
         when "000011001101" => index <= 5;
         when "000011001110" => index <= 5;
         when "000011001111" => index <= 4;
         when "000011010000" => index <= 7;
         when "000011010001" => index <= 5;
         when "000011010010" => index <= 6;
         when "000011010011" => index <= 5;
         when "000011010100" => index <= 6;
         when "000011010101" => index <= 5;
         when "000011010110" => index <= 5;
         when "000011010111" => index <= 4;
         when "000011011000" => index <= 6;
         when "000011011001" => index <= 5;
         when "000011011010" => index <= 5;
         when "000011011011" => index <= 4;
         when "000011011100" => index <= 5;
         when "000011011101" => index <= 5;
         when "000011011110" => index <= 5;
         when "000011011111" => index <= 4;
         when "000011100000" => index <= 7;
         when "000011100001" => index <= 6;
         when "000011100010" => index <= 6;
         when "000011100011" => index <= 5;
         when "000011100100" => index <= 6;
         when "000011100101" => index <= 5;
         when "000011100110" => index <= 5;
         when "000011100111" => index <= 4;
         when "000011101000" => index <= 6;
         when "000011101001" => index <= 5;
         when "000011101010" => index <= 5;
         when "000011101011" => index <= 5;
         when "000011101100" => index <= 6;
         when "000011101101" => index <= 5;
         when "000011101110" => index <= 5;
         when "000011101111" => index <= 4;
         when "000011110000" => index <= 6;
         when "000011110001" => index <= 5;
         when "000011110010" => index <= 6;
         when "000011110011" => index <= 5;
         when "000011110100" => index <= 6;
         when "000011110101" => index <= 5;
         when "000011110110" => index <= 5;
         when "000011110111" => index <= 5;
         when "000011111000" => index <= 6;
         when "000011111001" => index <= 5;
         when "000011111010" => index <= 5;
         when "000011111011" => index <= 5;
         when "000011111100" => index <= 6;
         when "000011111101" => index <= 5;
         when "000011111110" => index <= 5;
         when "000011111111" => index <= 4;
         when "000100000000" => index <= 9;
         when "000100000001" => index <= 5;
         when "000100000010" => index <= 6;
         when "000100000011" => index <= 4;
         when "000100000100" => index <= 6;
         when "000100000101" => index <= 4;
         when "000100000110" => index <= 5;
         when "000100000111" => index <= 4;
         when "000100001000" => index <= 6;
         when "000100001001" => index <= 5;
         when "000100001010" => index <= 5;
         when "000100001011" => index <= 4;
         when "000100001100" => index <= 5;
         when "000100001101" => index <= 4;
         when "000100001110" => index <= 4;
         when "000100001111" => index <= 4;
         when "000100010000" => index <= 7;
         when "000100010001" => index <= 5;
         when "000100010010" => index <= 5;
         when "000100010011" => index <= 4;
         when "000100010100" => index <= 6;
         when "000100010101" => index <= 4;
         when "000100010110" => index <= 5;
         when "000100010111" => index <= 4;
         when "000100011000" => index <= 6;
         when "000100011001" => index <= 5;
         when "000100011010" => index <= 5;
         when "000100011011" => index <= 4;
         when "000100011100" => index <= 5;
         when "000100011101" => index <= 4;
         when "000100011110" => index <= 5;
         when "000100011111" => index <= 4;
         when "000100100000" => index <= 8;
         when "000100100001" => index <= 5;
         when "000100100010" => index <= 6;
         when "000100100011" => index <= 4;
         when "000100100100" => index <= 6;
         when "000100100101" => index <= 5;
         when "000100100110" => index <= 5;
         when "000100100111" => index <= 4;
         when "000100101000" => index <= 6;
         when "000100101001" => index <= 5;
         when "000100101010" => index <= 5;
         when "000100101011" => index <= 4;
         when "000100101100" => index <= 6;
         when "000100101101" => index <= 5;
         when "000100101110" => index <= 5;
         when "000100101111" => index <= 4;
         when "000100110000" => index <= 7;
         when "000100110001" => index <= 5;
         when "000100110010" => index <= 6;
         when "000100110011" => index <= 5;
         when "000100110100" => index <= 6;
         when "000100110101" => index <= 5;
         when "000100110110" => index <= 5;
         when "000100110111" => index <= 4;
         when "000100111000" => index <= 6;
         when "000100111001" => index <= 5;
         when "000100111010" => index <= 5;
         when "000100111011" => index <= 4;
         when "000100111100" => index <= 5;
         when "000100111101" => index <= 5;
         when "000100111110" => index <= 5;
         when "000100111111" => index <= 4;
         when "000101000000" => index <= 8;
         when "000101000001" => index <= 6;
         when "000101000010" => index <= 6;
         when "000101000011" => index <= 5;
         when "000101000100" => index <= 6;
         when "000101000101" => index <= 5;
         when "000101000110" => index <= 5;
         when "000101000111" => index <= 4;
         when "000101001000" => index <= 7;
         when "000101001001" => index <= 5;
         when "000101001010" => index <= 6;
         when "000101001011" => index <= 5;
         when "000101001100" => index <= 6;
         when "000101001101" => index <= 5;
         when "000101001110" => index <= 5;
         when "000101001111" => index <= 4;
         when "000101010000" => index <= 7;
         when "000101010001" => index <= 6;
         when "000101010010" => index <= 6;
         when "000101010011" => index <= 5;
         when "000101010100" => index <= 6;
         when "000101010101" => index <= 5;
         when "000101010110" => index <= 5;
         when "000101010111" => index <= 4;
         when "000101011000" => index <= 6;
         when "000101011001" => index <= 5;
         when "000101011010" => index <= 5;
         when "000101011011" => index <= 5;
         when "000101011100" => index <= 6;
         when "000101011101" => index <= 5;
         when "000101011110" => index <= 5;
         when "000101011111" => index <= 4;
         when "000101100000" => index <= 7;
         when "000101100001" => index <= 6;
         when "000101100010" => index <= 6;
         when "000101100011" => index <= 5;
         when "000101100100" => index <= 6;
         when "000101100101" => index <= 5;
         when "000101100110" => index <= 5;
         when "000101100111" => index <= 5;
         when "000101101000" => index <= 6;
         when "000101101001" => index <= 5;
         when "000101101010" => index <= 6;
         when "000101101011" => index <= 5;
         when "000101101100" => index <= 6;
         when "000101101101" => index <= 5;
         when "000101101110" => index <= 5;
         when "000101101111" => index <= 5;
         when "000101110000" => index <= 7;
         when "000101110001" => index <= 6;
         when "000101110010" => index <= 6;
         when "000101110011" => index <= 5;
         when "000101110100" => index <= 6;
         when "000101110101" => index <= 5;
         when "000101110110" => index <= 5;
         when "000101110111" => index <= 5;
         when "000101111000" => index <= 6;
         when "000101111001" => index <= 5;
         when "000101111010" => index <= 6;
         when "000101111011" => index <= 5;
         when "000101111100" => index <= 6;
         when "000101111101" => index <= 5;
         when "000101111110" => index <= 5;
         when "000101111111" => index <= 5;
         when "000110000000" => index <= 8;
         when "000110000001" => index <= 6;
         when "000110000010" => index <= 6;
         when "000110000011" => index <= 5;
         when "000110000100" => index <= 7;
         when "000110000101" => index <= 5;
         when "000110000110" => index <= 6;
         when "000110000111" => index <= 5;
         when "000110001000" => index <= 7;
         when "000110001001" => index <= 6;
         when "000110001010" => index <= 6;
         when "000110001011" => index <= 5;
         when "000110001100" => index <= 6;
         when "000110001101" => index <= 5;
         when "000110001110" => index <= 5;
         when "000110001111" => index <= 4;
         when "000110010000" => index <= 7;
         when "000110010001" => index <= 6;
         when "000110010010" => index <= 6;
         when "000110010011" => index <= 5;
         when "000110010100" => index <= 6;
         when "000110010101" => index <= 5;
         when "000110010110" => index <= 5;
         when "000110010111" => index <= 5;
         when "000110011000" => index <= 6;
         when "000110011001" => index <= 5;
         when "000110011010" => index <= 6;
         when "000110011011" => index <= 5;
         when "000110011100" => index <= 6;
         when "000110011101" => index <= 5;
         when "000110011110" => index <= 5;
         when "000110011111" => index <= 5;
         when "000110100000" => index <= 8;
         when "000110100001" => index <= 6;
         when "000110100010" => index <= 6;
         when "000110100011" => index <= 5;
         when "000110100100" => index <= 6;
         when "000110100101" => index <= 5;
         when "000110100110" => index <= 6;
         when "000110100111" => index <= 5;
         when "000110101000" => index <= 7;
         when "000110101001" => index <= 6;
         when "000110101010" => index <= 6;
         when "000110101011" => index <= 5;
         when "000110101100" => index <= 6;
         when "000110101101" => index <= 5;
         when "000110101110" => index <= 5;
         when "000110101111" => index <= 5;
         when "000110110000" => index <= 7;
         when "000110110001" => index <= 6;
         when "000110110010" => index <= 6;
         when "000110110011" => index <= 5;
         when "000110110100" => index <= 6;
         when "000110110101" => index <= 5;
         when "000110110110" => index <= 6;
         when "000110110111" => index <= 5;
         when "000110111000" => index <= 6;
         when "000110111001" => index <= 6;
         when "000110111010" => index <= 6;
         when "000110111011" => index <= 5;
         when "000110111100" => index <= 6;
         when "000110111101" => index <= 5;
         when "000110111110" => index <= 5;
         when "000110111111" => index <= 5;
         when "000111000000" => index <= 8;
         when "000111000001" => index <= 6;
         when "000111000010" => index <= 6;
         when "000111000011" => index <= 5;
         when "000111000100" => index <= 7;
         when "000111000101" => index <= 6;
         when "000111000110" => index <= 6;
         when "000111000111" => index <= 5;
         when "000111001000" => index <= 7;
         when "000111001001" => index <= 6;
         when "000111001010" => index <= 6;
         when "000111001011" => index <= 5;
         when "000111001100" => index <= 6;
         when "000111001101" => index <= 5;
         when "000111001110" => index <= 6;
         when "000111001111" => index <= 5;
         when "000111010000" => index <= 7;
         when "000111010001" => index <= 6;
         when "000111010010" => index <= 6;
         when "000111010011" => index <= 5;
         when "000111010100" => index <= 6;
         when "000111010101" => index <= 6;
         when "000111010110" => index <= 6;
         when "000111010111" => index <= 5;
         when "000111011000" => index <= 7;
         when "000111011001" => index <= 6;
         when "000111011010" => index <= 6;
         when "000111011011" => index <= 5;
         when "000111011100" => index <= 6;
         when "000111011101" => index <= 5;
         when "000111011110" => index <= 5;
         when "000111011111" => index <= 5;
         when "000111100000" => index <= 8;
         when "000111100001" => index <= 6;
         when "000111100010" => index <= 6;
         when "000111100011" => index <= 6;
         when "000111100100" => index <= 7;
         when "000111100101" => index <= 6;
         when "000111100110" => index <= 6;
         when "000111100111" => index <= 5;
         when "000111101000" => index <= 7;
         when "000111101001" => index <= 6;
         when "000111101010" => index <= 6;
         when "000111101011" => index <= 5;
         when "000111101100" => index <= 6;
         when "000111101101" => index <= 5;
         when "000111101110" => index <= 6;
         when "000111101111" => index <= 5;
         when "000111110000" => index <= 7;
         when "000111110001" => index <= 6;
         when "000111110010" => index <= 6;
         when "000111110011" => index <= 5;
         when "000111110100" => index <= 6;
         when "000111110101" => index <= 6;
         when "000111110110" => index <= 6;
         when "000111110111" => index <= 5;
         when "000111111000" => index <= 6;
         when "000111111001" => index <= 6;
         when "000111111010" => index <= 6;
         when "000111111011" => index <= 5;
         when "000111111100" => index <= 6;
         when "000111111101" => index <= 5;
         when "000111111110" => index <= 6;
         when "000111111111" => index <= 5;
         when "001000000000" => index <= 10;
         when "001000000001" => index <= 6;
         when "001000000010" => index <= 6;
         when "001000000011" => index <= 4;
         when "001000000100" => index <= 6;
         when "001000000101" => index <= 5;
         when "001000000110" => index <= 5;
         when "001000000111" => index <= 4;
         when "001000001000" => index <= 7;
         when "001000001001" => index <= 5;
         when "001000001010" => index <= 5;
         when "001000001011" => index <= 4;
         when "001000001100" => index <= 6;
         when "001000001101" => index <= 4;
         when "001000001110" => index <= 5;
         when "001000001111" => index <= 4;
         when "001000010000" => index <= 8;
         when "001000010001" => index <= 5;
         when "001000010010" => index <= 6;
         when "001000010011" => index <= 4;
         when "001000010100" => index <= 6;
         when "001000010101" => index <= 5;
         when "001000010110" => index <= 5;
         when "001000010111" => index <= 4;
         when "001000011000" => index <= 6;
         when "001000011001" => index <= 5;
         when "001000011010" => index <= 5;
         when "001000011011" => index <= 4;
         when "001000011100" => index <= 6;
         when "001000011101" => index <= 5;
         when "001000011110" => index <= 5;
         when "001000011111" => index <= 4;
         when "001000100000" => index <= 8;
         when "001000100001" => index <= 6;
         when "001000100010" => index <= 6;
         when "001000100011" => index <= 5;
         when "001000100100" => index <= 6;
         when "001000100101" => index <= 5;
         when "001000100110" => index <= 5;
         when "001000100111" => index <= 4;
         when "001000101000" => index <= 7;
         when "001000101001" => index <= 5;
         when "001000101010" => index <= 6;
         when "001000101011" => index <= 5;
         when "001000101100" => index <= 6;
         when "001000101101" => index <= 5;
         when "001000101110" => index <= 5;
         when "001000101111" => index <= 4;
         when "001000110000" => index <= 7;
         when "001000110001" => index <= 6;
         when "001000110010" => index <= 6;
         when "001000110011" => index <= 5;
         when "001000110100" => index <= 6;
         when "001000110101" => index <= 5;
         when "001000110110" => index <= 5;
         when "001000110111" => index <= 4;
         when "001000111000" => index <= 6;
         when "001000111001" => index <= 5;
         when "001000111010" => index <= 5;
         when "001000111011" => index <= 5;
         when "001000111100" => index <= 6;
         when "001000111101" => index <= 5;
         when "001000111110" => index <= 5;
         when "001000111111" => index <= 4;
         when "001001000000" => index <= 8;
         when "001001000001" => index <= 6;
         when "001001000010" => index <= 6;
         when "001001000011" => index <= 5;
         when "001001000100" => index <= 7;
         when "001001000101" => index <= 5;
         when "001001000110" => index <= 6;
         when "001001000111" => index <= 5;
         when "001001001000" => index <= 7;
         when "001001001001" => index <= 6;
         when "001001001010" => index <= 6;
         when "001001001011" => index <= 5;
         when "001001001100" => index <= 6;
         when "001001001101" => index <= 5;
         when "001001001110" => index <= 5;
         when "001001001111" => index <= 4;
         when "001001010000" => index <= 7;
         when "001001010001" => index <= 6;
         when "001001010010" => index <= 6;
         when "001001010011" => index <= 5;
         when "001001010100" => index <= 6;
         when "001001010101" => index <= 5;
         when "001001010110" => index <= 5;
         when "001001010111" => index <= 5;
         when "001001011000" => index <= 6;
         when "001001011001" => index <= 5;
         when "001001011010" => index <= 6;
         when "001001011011" => index <= 5;
         when "001001011100" => index <= 6;
         when "001001011101" => index <= 5;
         when "001001011110" => index <= 5;
         when "001001011111" => index <= 5;
         when "001001100000" => index <= 8;
         when "001001100001" => index <= 6;
         when "001001100010" => index <= 6;
         when "001001100011" => index <= 5;
         when "001001100100" => index <= 6;
         when "001001100101" => index <= 5;
         when "001001100110" => index <= 6;
         when "001001100111" => index <= 5;
         when "001001101000" => index <= 7;
         when "001001101001" => index <= 6;
         when "001001101010" => index <= 6;
         when "001001101011" => index <= 5;
         when "001001101100" => index <= 6;
         when "001001101101" => index <= 5;
         when "001001101110" => index <= 5;
         when "001001101111" => index <= 5;
         when "001001110000" => index <= 7;
         when "001001110001" => index <= 6;
         when "001001110010" => index <= 6;
         when "001001110011" => index <= 5;
         when "001001110100" => index <= 6;
         when "001001110101" => index <= 5;
         when "001001110110" => index <= 6;
         when "001001110111" => index <= 5;
         when "001001111000" => index <= 6;
         when "001001111001" => index <= 6;
         when "001001111010" => index <= 6;
         when "001001111011" => index <= 5;
         when "001001111100" => index <= 6;
         when "001001111101" => index <= 5;
         when "001001111110" => index <= 5;
         when "001001111111" => index <= 5;
         when "001010000000" => index <= 9;
         when "001010000001" => index <= 6;
         when "001010000010" => index <= 7;
         when "001010000011" => index <= 5;
         when "001010000100" => index <= 7;
         when "001010000101" => index <= 6;
         when "001010000110" => index <= 6;
         when "001010000111" => index <= 5;
         when "001010001000" => index <= 7;
         when "001010001001" => index <= 6;
         when "001010001010" => index <= 6;
         when "001010001011" => index <= 5;
         when "001010001100" => index <= 6;
         when "001010001101" => index <= 5;
         when "001010001110" => index <= 5;
         when "001010001111" => index <= 5;
         when "001010010000" => index <= 8;
         when "001010010001" => index <= 6;
         when "001010010010" => index <= 6;
         when "001010010011" => index <= 5;
         when "001010010100" => index <= 6;
         when "001010010101" => index <= 5;
         when "001010010110" => index <= 6;
         when "001010010111" => index <= 5;
         when "001010011000" => index <= 7;
         when "001010011001" => index <= 6;
         when "001010011010" => index <= 6;
         when "001010011011" => index <= 5;
         when "001010011100" => index <= 6;
         when "001010011101" => index <= 5;
         when "001010011110" => index <= 5;
         when "001010011111" => index <= 5;
         when "001010100000" => index <= 8;
         when "001010100001" => index <= 6;
         when "001010100010" => index <= 6;
         when "001010100011" => index <= 5;
         when "001010100100" => index <= 7;
         when "001010100101" => index <= 6;
         when "001010100110" => index <= 6;
         when "001010100111" => index <= 5;
         when "001010101000" => index <= 7;
         when "001010101001" => index <= 6;
         when "001010101010" => index <= 6;
         when "001010101011" => index <= 5;
         when "001010101100" => index <= 6;
         when "001010101101" => index <= 5;
         when "001010101110" => index <= 6;
         when "001010101111" => index <= 5;
         when "001010110000" => index <= 7;
         when "001010110001" => index <= 6;
         when "001010110010" => index <= 6;
         when "001010110011" => index <= 5;
         when "001010110100" => index <= 6;
         when "001010110101" => index <= 6;
         when "001010110110" => index <= 6;
         when "001010110111" => index <= 5;
         when "001010111000" => index <= 7;
         when "001010111001" => index <= 6;
         when "001010111010" => index <= 6;
         when "001010111011" => index <= 5;
         when "001010111100" => index <= 6;
         when "001010111101" => index <= 5;
         when "001010111110" => index <= 5;
         when "001010111111" => index <= 5;
         when "001011000000" => index <= 8;
         when "001011000001" => index <= 6;
         when "001011000010" => index <= 7;
         when "001011000011" => index <= 6;
         when "001011000100" => index <= 7;
         when "001011000101" => index <= 6;
         when "001011000110" => index <= 6;
         when "001011000111" => index <= 5;
         when "001011001000" => index <= 7;
         when "001011001001" => index <= 6;
         when "001011001010" => index <= 6;
         when "001011001011" => index <= 5;
         when "001011001100" => index <= 6;
         when "001011001101" => index <= 6;
         when "001011001110" => index <= 6;
         when "001011001111" => index <= 5;
         when "001011010000" => index <= 8;
         when "001011010001" => index <= 6;
         when "001011010010" => index <= 6;
         when "001011010011" => index <= 6;
         when "001011010100" => index <= 7;
         when "001011010101" => index <= 6;
         when "001011010110" => index <= 6;
         when "001011010111" => index <= 5;
         when "001011011000" => index <= 7;
         when "001011011001" => index <= 6;
         when "001011011010" => index <= 6;
         when "001011011011" => index <= 5;
         when "001011011100" => index <= 6;
         when "001011011101" => index <= 5;
         when "001011011110" => index <= 6;
         when "001011011111" => index <= 5;
         when "001011100000" => index <= 8;
         when "001011100001" => index <= 6;
         when "001011100010" => index <= 7;
         when "001011100011" => index <= 6;
         when "001011100100" => index <= 7;
         when "001011100101" => index <= 6;
         when "001011100110" => index <= 6;
         when "001011100111" => index <= 5;
         when "001011101000" => index <= 7;
         when "001011101001" => index <= 6;
         when "001011101010" => index <= 6;
         when "001011101011" => index <= 5;
         when "001011101100" => index <= 6;
         when "001011101101" => index <= 6;
         when "001011101110" => index <= 6;
         when "001011101111" => index <= 5;
         when "001011110000" => index <= 7;
         when "001011110001" => index <= 6;
         when "001011110010" => index <= 6;
         when "001011110011" => index <= 6;
         when "001011110100" => index <= 6;
         when "001011110101" => index <= 6;
         when "001011110110" => index <= 6;
         when "001011110111" => index <= 5;
         when "001011111000" => index <= 7;
         when "001011111001" => index <= 6;
         when "001011111010" => index <= 6;
         when "001011111011" => index <= 5;
         when "001011111100" => index <= 6;
         when "001011111101" => index <= 6;
         when "001011111110" => index <= 6;
         when "001011111111" => index <= 5;
         when "001100000000" => index <= 10;
         when "001100000001" => index <= 7;
         when "001100000010" => index <= 7;
         when "001100000011" => index <= 6;
         when "001100000100" => index <= 7;
         when "001100000101" => index <= 6;
         when "001100000110" => index <= 6;
         when "001100000111" => index <= 5;
         when "001100001000" => index <= 8;
         when "001100001001" => index <= 6;
         when "001100001010" => index <= 6;
         when "001100001011" => index <= 5;
         when "001100001100" => index <= 6;
         when "001100001101" => index <= 5;
         when "001100001110" => index <= 6;
         when "001100001111" => index <= 5;
         when "001100010000" => index <= 8;
         when "001100010001" => index <= 6;
         when "001100010010" => index <= 6;
         when "001100010011" => index <= 5;
         when "001100010100" => index <= 7;
         when "001100010101" => index <= 6;
         when "001100010110" => index <= 6;
         when "001100010111" => index <= 5;
         when "001100011000" => index <= 7;
         when "001100011001" => index <= 6;
         when "001100011010" => index <= 6;
         when "001100011011" => index <= 5;
         when "001100011100" => index <= 6;
         when "001100011101" => index <= 5;
         when "001100011110" => index <= 6;
         when "001100011111" => index <= 5;
         when "001100100000" => index <= 8;
         when "001100100001" => index <= 6;
         when "001100100010" => index <= 7;
         when "001100100011" => index <= 6;
         when "001100100100" => index <= 7;
         when "001100100101" => index <= 6;
         when "001100100110" => index <= 6;
         when "001100100111" => index <= 5;
         when "001100101000" => index <= 7;
         when "001100101001" => index <= 6;
         when "001100101010" => index <= 6;
         when "001100101011" => index <= 5;
         when "001100101100" => index <= 6;
         when "001100101101" => index <= 6;
         when "001100101110" => index <= 6;
         when "001100101111" => index <= 5;
         when "001100110000" => index <= 8;
         when "001100110001" => index <= 6;
         when "001100110010" => index <= 6;
         when "001100110011" => index <= 6;
         when "001100110100" => index <= 7;
         when "001100110101" => index <= 6;
         when "001100110110" => index <= 6;
         when "001100110111" => index <= 5;
         when "001100111000" => index <= 7;
         when "001100111001" => index <= 6;
         when "001100111010" => index <= 6;
         when "001100111011" => index <= 5;
         when "001100111100" => index <= 6;
         when "001100111101" => index <= 5;
         when "001100111110" => index <= 6;
         when "001100111111" => index <= 5;
         when "001101000000" => index <= 9;
         when "001101000001" => index <= 7;
         when "001101000010" => index <= 7;
         when "001101000011" => index <= 6;
         when "001101000100" => index <= 7;
         when "001101000101" => index <= 6;
         when "001101000110" => index <= 6;
         when "001101000111" => index <= 5;
         when "001101001000" => index <= 8;
         when "001101001001" => index <= 6;
         when "001101001010" => index <= 6;
         when "001101001011" => index <= 6;
         when "001101001100" => index <= 7;
         when "001101001101" => index <= 6;
         when "001101001110" => index <= 6;
         when "001101001111" => index <= 5;
         when "001101010000" => index <= 8;
         when "001101010001" => index <= 6;
         when "001101010010" => index <= 7;
         when "001101010011" => index <= 6;
         when "001101010100" => index <= 7;
         when "001101010101" => index <= 6;
         when "001101010110" => index <= 6;
         when "001101010111" => index <= 5;
         when "001101011000" => index <= 7;
         when "001101011001" => index <= 6;
         when "001101011010" => index <= 6;
         when "001101011011" => index <= 5;
         when "001101011100" => index <= 6;
         when "001101011101" => index <= 6;
         when "001101011110" => index <= 6;
         when "001101011111" => index <= 5;
         when "001101100000" => index <= 8;
         when "001101100001" => index <= 7;
         when "001101100010" => index <= 7;
         when "001101100011" => index <= 6;
         when "001101100100" => index <= 7;
         when "001101100101" => index <= 6;
         when "001101100110" => index <= 6;
         when "001101100111" => index <= 5;
         when "001101101000" => index <= 7;
         when "001101101001" => index <= 6;
         when "001101101010" => index <= 6;
         when "001101101011" => index <= 6;
         when "001101101100" => index <= 6;
         when "001101101101" => index <= 6;
         when "001101101110" => index <= 6;
         when "001101101111" => index <= 5;
         when "001101110000" => index <= 7;
         when "001101110001" => index <= 6;
         when "001101110010" => index <= 6;
         when "001101110011" => index <= 6;
         when "001101110100" => index <= 7;
         when "001101110101" => index <= 6;
         when "001101110110" => index <= 6;
         when "001101110111" => index <= 5;
         when "001101111000" => index <= 7;
         when "001101111001" => index <= 6;
         when "001101111010" => index <= 6;
         when "001101111011" => index <= 6;
         when "001101111100" => index <= 6;
         when "001101111101" => index <= 6;
         when "001101111110" => index <= 6;
         when "001101111111" => index <= 5;
         when "001110000000" => index <= 9;
         when "001110000001" => index <= 7;
         when "001110000010" => index <= 7;
         when "001110000011" => index <= 6;
         when "001110000100" => index <= 8;
         when "001110000101" => index <= 6;
         when "001110000110" => index <= 6;
         when "001110000111" => index <= 6;
         when "001110001000" => index <= 8;
         when "001110001001" => index <= 6;
         when "001110001010" => index <= 7;
         when "001110001011" => index <= 6;
         when "001110001100" => index <= 7;
         when "001110001101" => index <= 6;
         when "001110001110" => index <= 6;
         when "001110001111" => index <= 5;
         when "001110010000" => index <= 8;
         when "001110010001" => index <= 7;
         when "001110010010" => index <= 7;
         when "001110010011" => index <= 6;
         when "001110010100" => index <= 7;
         when "001110010101" => index <= 6;
         when "001110010110" => index <= 6;
         when "001110010111" => index <= 5;
         when "001110011000" => index <= 7;
         when "001110011001" => index <= 6;
         when "001110011010" => index <= 6;
         when "001110011011" => index <= 6;
         when "001110011100" => index <= 6;
         when "001110011101" => index <= 6;
         when "001110011110" => index <= 6;
         when "001110011111" => index <= 5;
         when "001110100000" => index <= 8;
         when "001110100001" => index <= 7;
         when "001110100010" => index <= 7;
         when "001110100011" => index <= 6;
         when "001110100100" => index <= 7;
         when "001110100101" => index <= 6;
         when "001110100110" => index <= 6;
         when "001110100111" => index <= 6;
         when "001110101000" => index <= 7;
         when "001110101001" => index <= 6;
         when "001110101010" => index <= 6;
         when "001110101011" => index <= 6;
         when "001110101100" => index <= 7;
         when "001110101101" => index <= 6;
         when "001110101110" => index <= 6;
         when "001110101111" => index <= 5;
         when "001110110000" => index <= 8;
         when "001110110001" => index <= 6;
         when "001110110010" => index <= 7;
         when "001110110011" => index <= 6;
         when "001110110100" => index <= 7;
         when "001110110101" => index <= 6;
         when "001110110110" => index <= 6;
         when "001110110111" => index <= 6;
         when "001110111000" => index <= 7;
         when "001110111001" => index <= 6;
         when "001110111010" => index <= 6;
         when "001110111011" => index <= 6;
         when "001110111100" => index <= 6;
         when "001110111101" => index <= 6;
         when "001110111110" => index <= 6;
         when "001110111111" => index <= 5;
         when "001111000000" => index <= 8;
         when "001111000001" => index <= 7;
         when "001111000010" => index <= 7;
         when "001111000011" => index <= 6;
         when "001111000100" => index <= 7;
         when "001111000101" => index <= 6;
         when "001111000110" => index <= 6;
         when "001111000111" => index <= 6;
         when "001111001000" => index <= 8;
         when "001111001001" => index <= 6;
         when "001111001010" => index <= 7;
         when "001111001011" => index <= 6;
         when "001111001100" => index <= 7;
         when "001111001101" => index <= 6;
         when "001111001110" => index <= 6;
         when "001111001111" => index <= 6;
         when "001111010000" => index <= 8;
         when "001111010001" => index <= 7;
         when "001111010010" => index <= 7;
         when "001111010011" => index <= 6;
         when "001111010100" => index <= 7;
         when "001111010101" => index <= 6;
         when "001111010110" => index <= 6;
         when "001111010111" => index <= 6;
         when "001111011000" => index <= 7;
         when "001111011001" => index <= 6;
         when "001111011010" => index <= 6;
         when "001111011011" => index <= 6;
         when "001111011100" => index <= 7;
         when "001111011101" => index <= 6;
         when "001111011110" => index <= 6;
         when "001111011111" => index <= 5;
         when "001111100000" => index <= 8;
         when "001111100001" => index <= 7;
         when "001111100010" => index <= 7;
         when "001111100011" => index <= 6;
         when "001111100100" => index <= 7;
         when "001111100101" => index <= 6;
         when "001111100110" => index <= 6;
         when "001111100111" => index <= 6;
         when "001111101000" => index <= 7;
         when "001111101001" => index <= 6;
         when "001111101010" => index <= 7;
         when "001111101011" => index <= 6;
         when "001111101100" => index <= 7;
         when "001111101101" => index <= 6;
         when "001111101110" => index <= 6;
         when "001111101111" => index <= 6;
         when "001111110000" => index <= 8;
         when "001111110001" => index <= 7;
         when "001111110010" => index <= 7;
         when "001111110011" => index <= 6;
         when "001111110100" => index <= 7;
         when "001111110101" => index <= 6;
         when "001111110110" => index <= 6;
         when "001111110111" => index <= 6;
         when "001111111000" => index <= 7;
         when "001111111001" => index <= 6;
         when "001111111010" => index <= 6;
         when "001111111011" => index <= 6;
         when "001111111100" => index <= 6;
         when "001111111101" => index <= 6;
         when "001111111110" => index <= 6;
         when "001111111111" => index <= 6;
         when "010000000000" => index <= 11;
         when "010000000001" => index <= 6;
         when "010000000010" => index <= 6;
         when "010000000011" => index <= 5;
         when "010000000100" => index <= 7;
         when "010000000101" => index <= 5;
         when "010000000110" => index <= 5;
         when "010000000111" => index <= 4;
         when "010000001000" => index <= 8;
         when "010000001001" => index <= 5;
         when "010000001010" => index <= 6;
         when "010000001011" => index <= 4;
         when "010000001100" => index <= 6;
         when "010000001101" => index <= 5;
         when "010000001110" => index <= 5;
         when "010000001111" => index <= 4;
         when "010000010000" => index <= 8;
         when "010000010001" => index <= 6;
         when "010000010010" => index <= 6;
         when "010000010011" => index <= 5;
         when "010000010100" => index <= 6;
         when "010000010101" => index <= 5;
         when "010000010110" => index <= 5;
         when "010000010111" => index <= 4;
         when "010000011000" => index <= 7;
         when "010000011001" => index <= 5;
         when "010000011010" => index <= 6;
         when "010000011011" => index <= 5;
         when "010000011100" => index <= 6;
         when "010000011101" => index <= 5;
         when "010000011110" => index <= 5;
         when "010000011111" => index <= 4;
         when "010000100000" => index <= 8;
         when "010000100001" => index <= 6;
         when "010000100010" => index <= 6;
         when "010000100011" => index <= 5;
         when "010000100100" => index <= 7;
         when "010000100101" => index <= 5;
         when "010000100110" => index <= 6;
         when "010000100111" => index <= 5;
         when "010000101000" => index <= 7;
         when "010000101001" => index <= 6;
         when "010000101010" => index <= 6;
         when "010000101011" => index <= 5;
         when "010000101100" => index <= 6;
         when "010000101101" => index <= 5;
         when "010000101110" => index <= 5;
         when "010000101111" => index <= 4;
         when "010000110000" => index <= 7;
         when "010000110001" => index <= 6;
         when "010000110010" => index <= 6;
         when "010000110011" => index <= 5;
         when "010000110100" => index <= 6;
         when "010000110101" => index <= 5;
         when "010000110110" => index <= 5;
         when "010000110111" => index <= 5;
         when "010000111000" => index <= 6;
         when "010000111001" => index <= 5;
         when "010000111010" => index <= 6;
         when "010000111011" => index <= 5;
         when "010000111100" => index <= 6;
         when "010000111101" => index <= 5;
         when "010000111110" => index <= 5;
         when "010000111111" => index <= 5;
         when "010001000000" => index <= 9;
         when "010001000001" => index <= 6;
         when "010001000010" => index <= 7;
         when "010001000011" => index <= 5;
         when "010001000100" => index <= 7;
         when "010001000101" => index <= 6;
         when "010001000110" => index <= 6;
         when "010001000111" => index <= 5;
         when "010001001000" => index <= 7;
         when "010001001001" => index <= 6;
         when "010001001010" => index <= 6;
         when "010001001011" => index <= 5;
         when "010001001100" => index <= 6;
         when "010001001101" => index <= 5;
         when "010001001110" => index <= 5;
         when "010001001111" => index <= 5;
         when "010001010000" => index <= 8;
         when "010001010001" => index <= 6;
         when "010001010010" => index <= 6;
         when "010001010011" => index <= 5;
         when "010001010100" => index <= 6;
         when "010001010101" => index <= 5;
         when "010001010110" => index <= 6;
         when "010001010111" => index <= 5;
         when "010001011000" => index <= 7;
         when "010001011001" => index <= 6;
         when "010001011010" => index <= 6;
         when "010001011011" => index <= 5;
         when "010001011100" => index <= 6;
         when "010001011101" => index <= 5;
         when "010001011110" => index <= 5;
         when "010001011111" => index <= 5;
         when "010001100000" => index <= 8;
         when "010001100001" => index <= 6;
         when "010001100010" => index <= 6;
         when "010001100011" => index <= 5;
         when "010001100100" => index <= 7;
         when "010001100101" => index <= 6;
         when "010001100110" => index <= 6;
         when "010001100111" => index <= 5;
         when "010001101000" => index <= 7;
         when "010001101001" => index <= 6;
         when "010001101010" => index <= 6;
         when "010001101011" => index <= 5;
         when "010001101100" => index <= 6;
         when "010001101101" => index <= 5;
         when "010001101110" => index <= 6;
         when "010001101111" => index <= 5;
         when "010001110000" => index <= 7;
         when "010001110001" => index <= 6;
         when "010001110010" => index <= 6;
         when "010001110011" => index <= 5;
         when "010001110100" => index <= 6;
         when "010001110101" => index <= 6;
         when "010001110110" => index <= 6;
         when "010001110111" => index <= 5;
         when "010001111000" => index <= 7;
         when "010001111001" => index <= 6;
         when "010001111010" => index <= 6;
         when "010001111011" => index <= 5;
         when "010001111100" => index <= 6;
         when "010001111101" => index <= 5;
         when "010001111110" => index <= 5;
         when "010001111111" => index <= 5;
         when "010010000000" => index <= 10;
         when "010010000001" => index <= 7;
         when "010010000010" => index <= 7;
         when "010010000011" => index <= 6;
         when "010010000100" => index <= 7;
         when "010010000101" => index <= 6;
         when "010010000110" => index <= 6;
         when "010010000111" => index <= 5;
         when "010010001000" => index <= 8;
         when "010010001001" => index <= 6;
         when "010010001010" => index <= 6;
         when "010010001011" => index <= 5;
         when "010010001100" => index <= 6;
         when "010010001101" => index <= 5;
         when "010010001110" => index <= 6;
         when "010010001111" => index <= 5;
         when "010010010000" => index <= 8;
         when "010010010001" => index <= 6;
         when "010010010010" => index <= 6;
         when "010010010011" => index <= 5;
         when "010010010100" => index <= 7;
         when "010010010101" => index <= 6;
         when "010010010110" => index <= 6;
         when "010010010111" => index <= 5;
         when "010010011000" => index <= 7;
         when "010010011001" => index <= 6;
         when "010010011010" => index <= 6;
         when "010010011011" => index <= 5;
         when "010010011100" => index <= 6;
         when "010010011101" => index <= 5;
         when "010010011110" => index <= 6;
         when "010010011111" => index <= 5;
         when "010010100000" => index <= 8;
         when "010010100001" => index <= 6;
         when "010010100010" => index <= 7;
         when "010010100011" => index <= 6;
         when "010010100100" => index <= 7;
         when "010010100101" => index <= 6;
         when "010010100110" => index <= 6;
         when "010010100111" => index <= 5;
         when "010010101000" => index <= 7;
         when "010010101001" => index <= 6;
         when "010010101010" => index <= 6;
         when "010010101011" => index <= 5;
         when "010010101100" => index <= 6;
         when "010010101101" => index <= 6;
         when "010010101110" => index <= 6;
         when "010010101111" => index <= 5;
         when "010010110000" => index <= 8;
         when "010010110001" => index <= 6;
         when "010010110010" => index <= 6;
         when "010010110011" => index <= 6;
         when "010010110100" => index <= 7;
         when "010010110101" => index <= 6;
         when "010010110110" => index <= 6;
         when "010010110111" => index <= 5;
         when "010010111000" => index <= 7;
         when "010010111001" => index <= 6;
         when "010010111010" => index <= 6;
         when "010010111011" => index <= 5;
         when "010010111100" => index <= 6;
         when "010010111101" => index <= 5;
         when "010010111110" => index <= 6;
         when "010010111111" => index <= 5;
         when "010011000000" => index <= 9;
         when "010011000001" => index <= 7;
         when "010011000010" => index <= 7;
         when "010011000011" => index <= 6;
         when "010011000100" => index <= 7;
         when "010011000101" => index <= 6;
         when "010011000110" => index <= 6;
         when "010011000111" => index <= 5;
         when "010011001000" => index <= 8;
         when "010011001001" => index <= 6;
         when "010011001010" => index <= 6;
         when "010011001011" => index <= 6;
         when "010011001100" => index <= 7;
         when "010011001101" => index <= 6;
         when "010011001110" => index <= 6;
         when "010011001111" => index <= 5;
         when "010011010000" => index <= 8;
         when "010011010001" => index <= 6;
         when "010011010010" => index <= 7;
         when "010011010011" => index <= 6;
         when "010011010100" => index <= 7;
         when "010011010101" => index <= 6;
         when "010011010110" => index <= 6;
         when "010011010111" => index <= 5;
         when "010011011000" => index <= 7;
         when "010011011001" => index <= 6;
         when "010011011010" => index <= 6;
         when "010011011011" => index <= 5;
         when "010011011100" => index <= 6;
         when "010011011101" => index <= 6;
         when "010011011110" => index <= 6;
         when "010011011111" => index <= 5;
         when "010011100000" => index <= 8;
         when "010011100001" => index <= 7;
         when "010011100010" => index <= 7;
         when "010011100011" => index <= 6;
         when "010011100100" => index <= 7;
         when "010011100101" => index <= 6;
         when "010011100110" => index <= 6;
         when "010011100111" => index <= 5;
         when "010011101000" => index <= 7;
         when "010011101001" => index <= 6;
         when "010011101010" => index <= 6;
         when "010011101011" => index <= 6;
         when "010011101100" => index <= 6;
         when "010011101101" => index <= 6;
         when "010011101110" => index <= 6;
         when "010011101111" => index <= 5;
         when "010011110000" => index <= 7;
         when "010011110001" => index <= 6;
         when "010011110010" => index <= 6;
         when "010011110011" => index <= 6;
         when "010011110100" => index <= 7;
         when "010011110101" => index <= 6;
         when "010011110110" => index <= 6;
         when "010011110111" => index <= 5;
         when "010011111000" => index <= 7;
         when "010011111001" => index <= 6;
         when "010011111010" => index <= 6;
         when "010011111011" => index <= 6;
         when "010011111100" => index <= 6;
         when "010011111101" => index <= 6;
         when "010011111110" => index <= 6;
         when "010011111111" => index <= 5;
         when "010100000000" => index <= 10;
         when "010100000001" => index <= 7;
         when "010100000010" => index <= 7;
         when "010100000011" => index <= 6;
         when "010100000100" => index <= 8;
         when "010100000101" => index <= 6;
         when "010100000110" => index <= 6;
         when "010100000111" => index <= 5;
         when "010100001000" => index <= 8;
         when "010100001001" => index <= 6;
         when "010100001010" => index <= 6;
         when "010100001011" => index <= 5;
         when "010100001100" => index <= 7;
         when "010100001101" => index <= 6;
         when "010100001110" => index <= 6;
         when "010100001111" => index <= 5;
         when "010100010000" => index <= 8;
         when "010100010001" => index <= 6;
         when "010100010010" => index <= 7;
         when "010100010011" => index <= 6;
         when "010100010100" => index <= 7;
         when "010100010101" => index <= 6;
         when "010100010110" => index <= 6;
         when "010100010111" => index <= 5;
         when "010100011000" => index <= 7;
         when "010100011001" => index <= 6;
         when "010100011010" => index <= 6;
         when "010100011011" => index <= 5;
         when "010100011100" => index <= 6;
         when "010100011101" => index <= 6;
         when "010100011110" => index <= 6;
         when "010100011111" => index <= 5;
         when "010100100000" => index <= 9;
         when "010100100001" => index <= 7;
         when "010100100010" => index <= 7;
         when "010100100011" => index <= 6;
         when "010100100100" => index <= 7;
         when "010100100101" => index <= 6;
         when "010100100110" => index <= 6;
         when "010100100111" => index <= 5;
         when "010100101000" => index <= 8;
         when "010100101001" => index <= 6;
         when "010100101010" => index <= 6;
         when "010100101011" => index <= 6;
         when "010100101100" => index <= 7;
         when "010100101101" => index <= 6;
         when "010100101110" => index <= 6;
         when "010100101111" => index <= 5;
         when "010100110000" => index <= 8;
         when "010100110001" => index <= 6;
         when "010100110010" => index <= 7;
         when "010100110011" => index <= 6;
         when "010100110100" => index <= 7;
         when "010100110101" => index <= 6;
         when "010100110110" => index <= 6;
         when "010100110111" => index <= 5;
         when "010100111000" => index <= 7;
         when "010100111001" => index <= 6;
         when "010100111010" => index <= 6;
         when "010100111011" => index <= 5;
         when "010100111100" => index <= 6;
         when "010100111101" => index <= 6;
         when "010100111110" => index <= 6;
         when "010100111111" => index <= 5;
         when "010101000000" => index <= 9;
         when "010101000001" => index <= 7;
         when "010101000010" => index <= 7;
         when "010101000011" => index <= 6;
         when "010101000100" => index <= 8;
         when "010101000101" => index <= 6;
         when "010101000110" => index <= 6;
         when "010101000111" => index <= 6;
         when "010101001000" => index <= 8;
         when "010101001001" => index <= 6;
         when "010101001010" => index <= 7;
         when "010101001011" => index <= 6;
         when "010101001100" => index <= 7;
         when "010101001101" => index <= 6;
         when "010101001110" => index <= 6;
         when "010101001111" => index <= 5;
         when "010101010000" => index <= 8;
         when "010101010001" => index <= 7;
         when "010101010010" => index <= 7;
         when "010101010011" => index <= 6;
         when "010101010100" => index <= 7;
         when "010101010101" => index <= 6;
         when "010101010110" => index <= 6;
         when "010101010111" => index <= 5;
         when "010101011000" => index <= 7;
         when "010101011001" => index <= 6;
         when "010101011010" => index <= 6;
         when "010101011011" => index <= 6;
         when "010101011100" => index <= 6;
         when "010101011101" => index <= 6;
         when "010101011110" => index <= 6;
         when "010101011111" => index <= 5;
         when "010101100000" => index <= 8;
         when "010101100001" => index <= 7;
         when "010101100010" => index <= 7;
         when "010101100011" => index <= 6;
         when "010101100100" => index <= 7;
         when "010101100101" => index <= 6;
         when "010101100110" => index <= 6;
         when "010101100111" => index <= 6;
         when "010101101000" => index <= 7;
         when "010101101001" => index <= 6;
         when "010101101010" => index <= 6;
         when "010101101011" => index <= 6;
         when "010101101100" => index <= 7;
         when "010101101101" => index <= 6;
         when "010101101110" => index <= 6;
         when "010101101111" => index <= 5;
         when "010101110000" => index <= 8;
         when "010101110001" => index <= 6;
         when "010101110010" => index <= 7;
         when "010101110011" => index <= 6;
         when "010101110100" => index <= 7;
         when "010101110101" => index <= 6;
         when "010101110110" => index <= 6;
         when "010101110111" => index <= 6;
         when "010101111000" => index <= 7;
         when "010101111001" => index <= 6;
         when "010101111010" => index <= 6;
         when "010101111011" => index <= 6;
         when "010101111100" => index <= 6;
         when "010101111101" => index <= 6;
         when "010101111110" => index <= 6;
         when "010101111111" => index <= 5;
         when "010110000000" => index <= 9;
         when "010110000001" => index <= 7;
         when "010110000010" => index <= 8;
         when "010110000011" => index <= 6;
         when "010110000100" => index <= 8;
         when "010110000101" => index <= 6;
         when "010110000110" => index <= 7;
         when "010110000111" => index <= 6;
         when "010110001000" => index <= 8;
         when "010110001001" => index <= 7;
         when "010110001010" => index <= 7;
         when "010110001011" => index <= 6;
         when "010110001100" => index <= 7;
         when "010110001101" => index <= 6;
         when "010110001110" => index <= 6;
         when "010110001111" => index <= 5;
         when "010110010000" => index <= 8;
         when "010110010001" => index <= 7;
         when "010110010010" => index <= 7;
         when "010110010011" => index <= 6;
         when "010110010100" => index <= 7;
         when "010110010101" => index <= 6;
         when "010110010110" => index <= 6;
         when "010110010111" => index <= 6;
         when "010110011000" => index <= 7;
         when "010110011001" => index <= 6;
         when "010110011010" => index <= 6;
         when "010110011011" => index <= 6;
         when "010110011100" => index <= 7;
         when "010110011101" => index <= 6;
         when "010110011110" => index <= 6;
         when "010110011111" => index <= 5;
         when "010110100000" => index <= 8;
         when "010110100001" => index <= 7;
         when "010110100010" => index <= 7;
         when "010110100011" => index <= 6;
         when "010110100100" => index <= 7;
         when "010110100101" => index <= 6;
         when "010110100110" => index <= 6;
         when "010110100111" => index <= 6;
         when "010110101000" => index <= 8;
         when "010110101001" => index <= 6;
         when "010110101010" => index <= 7;
         when "010110101011" => index <= 6;
         when "010110101100" => index <= 7;
         when "010110101101" => index <= 6;
         when "010110101110" => index <= 6;
         when "010110101111" => index <= 6;
         when "010110110000" => index <= 8;
         when "010110110001" => index <= 7;
         when "010110110010" => index <= 7;
         when "010110110011" => index <= 6;
         when "010110110100" => index <= 7;
         when "010110110101" => index <= 6;
         when "010110110110" => index <= 6;
         when "010110110111" => index <= 6;
         when "010110111000" => index <= 7;
         when "010110111001" => index <= 6;
         when "010110111010" => index <= 6;
         when "010110111011" => index <= 6;
         when "010110111100" => index <= 7;
         when "010110111101" => index <= 6;
         when "010110111110" => index <= 6;
         when "010110111111" => index <= 5;
         when "010111000000" => index <= 9;
         when "010111000001" => index <= 7;
         when "010111000010" => index <= 7;
         when "010111000011" => index <= 6;
         when "010111000100" => index <= 8;
         when "010111000101" => index <= 6;
         when "010111000110" => index <= 7;
         when "010111000111" => index <= 6;
         when "010111001000" => index <= 8;
         when "010111001001" => index <= 7;
         when "010111001010" => index <= 7;
         when "010111001011" => index <= 6;
         when "010111001100" => index <= 7;
         when "010111001101" => index <= 6;
         when "010111001110" => index <= 6;
         when "010111001111" => index <= 6;
         when "010111010000" => index <= 8;
         when "010111010001" => index <= 7;
         when "010111010010" => index <= 7;
         when "010111010011" => index <= 6;
         when "010111010100" => index <= 7;
         when "010111010101" => index <= 6;
         when "010111010110" => index <= 6;
         when "010111010111" => index <= 6;
         when "010111011000" => index <= 7;
         when "010111011001" => index <= 6;
         when "010111011010" => index <= 7;
         when "010111011011" => index <= 6;
         when "010111011100" => index <= 7;
         when "010111011101" => index <= 6;
         when "010111011110" => index <= 6;
         when "010111011111" => index <= 6;
         when "010111100000" => index <= 8;
         when "010111100001" => index <= 7;
         when "010111100010" => index <= 7;
         when "010111100011" => index <= 6;
         when "010111100100" => index <= 7;
         when "010111100101" => index <= 6;
         when "010111100110" => index <= 7;
         when "010111100111" => index <= 6;
         when "010111101000" => index <= 8;
         when "010111101001" => index <= 7;
         when "010111101010" => index <= 7;
         when "010111101011" => index <= 6;
         when "010111101100" => index <= 7;
         when "010111101101" => index <= 6;
         when "010111101110" => index <= 6;
         when "010111101111" => index <= 6;
         when "010111110000" => index <= 8;
         when "010111110001" => index <= 7;
         when "010111110010" => index <= 7;
         when "010111110011" => index <= 6;
         when "010111110100" => index <= 7;
         when "010111110101" => index <= 6;
         when "010111110110" => index <= 6;
         when "010111110111" => index <= 6;
         when "010111111000" => index <= 7;
         when "010111111001" => index <= 6;
         when "010111111010" => index <= 6;
         when "010111111011" => index <= 6;
         when "010111111100" => index <= 7;
         when "010111111101" => index <= 6;
         when "010111111110" => index <= 6;
         when "010111111111" => index <= 6;
         when "011000000000" => index <= 10;
         when "011000000001" => index <= 7;
         when "011000000010" => index <= 8;
         when "011000000011" => index <= 6;
         when "011000000100" => index <= 8;
         when "011000000101" => index <= 6;
         when "011000000110" => index <= 6;
         when "011000000111" => index <= 5;
         when "011000001000" => index <= 8;
         when "011000001001" => index <= 6;
         when "011000001010" => index <= 7;
         when "011000001011" => index <= 6;
         when "011000001100" => index <= 7;
         when "011000001101" => index <= 6;
         when "011000001110" => index <= 6;
         when "011000001111" => index <= 5;
         when "011000010000" => index <= 9;
         when "011000010001" => index <= 7;
         when "011000010010" => index <= 7;
         when "011000010011" => index <= 6;
         when "011000010100" => index <= 7;
         when "011000010101" => index <= 6;
         when "011000010110" => index <= 6;
         when "011000010111" => index <= 5;
         when "011000011000" => index <= 8;
         when "011000011001" => index <= 6;
         when "011000011010" => index <= 6;
         when "011000011011" => index <= 6;
         when "011000011100" => index <= 7;
         when "011000011101" => index <= 6;
         when "011000011110" => index <= 6;
         when "011000011111" => index <= 5;
         when "011000100000" => index <= 9;
         when "011000100001" => index <= 7;
         when "011000100010" => index <= 7;
         when "011000100011" => index <= 6;
         when "011000100100" => index <= 8;
         when "011000100101" => index <= 6;
         when "011000100110" => index <= 6;
         when "011000100111" => index <= 6;
         when "011000101000" => index <= 8;
         when "011000101001" => index <= 6;
         when "011000101010" => index <= 7;
         when "011000101011" => index <= 6;
         when "011000101100" => index <= 7;
         when "011000101101" => index <= 6;
         when "011000101110" => index <= 6;
         when "011000101111" => index <= 5;
         when "011000110000" => index <= 8;
         when "011000110001" => index <= 7;
         when "011000110010" => index <= 7;
         when "011000110011" => index <= 6;
         when "011000110100" => index <= 7;
         when "011000110101" => index <= 6;
         when "011000110110" => index <= 6;
         when "011000110111" => index <= 5;
         when "011000111000" => index <= 7;
         when "011000111001" => index <= 6;
         when "011000111010" => index <= 6;
         when "011000111011" => index <= 6;
         when "011000111100" => index <= 6;
         when "011000111101" => index <= 6;
         when "011000111110" => index <= 6;
         when "011000111111" => index <= 5;
         when "011001000000" => index <= 9;
         when "011001000001" => index <= 7;
         when "011001000010" => index <= 8;
         when "011001000011" => index <= 6;
         when "011001000100" => index <= 8;
         when "011001000101" => index <= 6;
         when "011001000110" => index <= 7;
         when "011001000111" => index <= 6;
         when "011001001000" => index <= 8;
         when "011001001001" => index <= 7;
         when "011001001010" => index <= 7;
         when "011001001011" => index <= 6;
         when "011001001100" => index <= 7;
         when "011001001101" => index <= 6;
         when "011001001110" => index <= 6;
         when "011001001111" => index <= 5;
         when "011001010000" => index <= 8;
         when "011001010001" => index <= 7;
         when "011001010010" => index <= 7;
         when "011001010011" => index <= 6;
         when "011001010100" => index <= 7;
         when "011001010101" => index <= 6;
         when "011001010110" => index <= 6;
         when "011001010111" => index <= 6;
         when "011001011000" => index <= 7;
         when "011001011001" => index <= 6;
         when "011001011010" => index <= 6;
         when "011001011011" => index <= 6;
         when "011001011100" => index <= 7;
         when "011001011101" => index <= 6;
         when "011001011110" => index <= 6;
         when "011001011111" => index <= 5;
         when "011001100000" => index <= 8;
         when "011001100001" => index <= 7;
         when "011001100010" => index <= 7;
         when "011001100011" => index <= 6;
         when "011001100100" => index <= 7;
         when "011001100101" => index <= 6;
         when "011001100110" => index <= 6;
         when "011001100111" => index <= 6;
         when "011001101000" => index <= 8;
         when "011001101001" => index <= 6;
         when "011001101010" => index <= 7;
         when "011001101011" => index <= 6;
         when "011001101100" => index <= 7;
         when "011001101101" => index <= 6;
         when "011001101110" => index <= 6;
         when "011001101111" => index <= 6;
         when "011001110000" => index <= 8;
         when "011001110001" => index <= 7;
         when "011001110010" => index <= 7;
         when "011001110011" => index <= 6;
         when "011001110100" => index <= 7;
         when "011001110101" => index <= 6;
         when "011001110110" => index <= 6;
         when "011001110111" => index <= 6;
         when "011001111000" => index <= 7;
         when "011001111001" => index <= 6;
         when "011001111010" => index <= 6;
         when "011001111011" => index <= 6;
         when "011001111100" => index <= 7;
         when "011001111101" => index <= 6;
         when "011001111110" => index <= 6;
         when "011001111111" => index <= 5;
         when "011010000000" => index <= 10;
         when "011010000001" => index <= 8;
         when "011010000010" => index <= 8;
         when "011010000011" => index <= 6;
         when "011010000100" => index <= 8;
         when "011010000101" => index <= 7;
         when "011010000110" => index <= 7;
         when "011010000111" => index <= 6;
         when "011010001000" => index <= 8;
         when "011010001001" => index <= 7;
         when "011010001010" => index <= 7;
         when "011010001011" => index <= 6;
         when "011010001100" => index <= 7;
         when "011010001101" => index <= 6;
         when "011010001110" => index <= 6;
         when "011010001111" => index <= 6;
         when "011010010000" => index <= 8;
         when "011010010001" => index <= 7;
         when "011010010010" => index <= 7;
         when "011010010011" => index <= 6;
         when "011010010100" => index <= 7;
         when "011010010101" => index <= 6;
         when "011010010110" => index <= 6;
         when "011010010111" => index <= 6;
         when "011010011000" => index <= 8;
         when "011010011001" => index <= 6;
         when "011010011010" => index <= 7;
         when "011010011011" => index <= 6;
         when "011010011100" => index <= 7;
         when "011010011101" => index <= 6;
         when "011010011110" => index <= 6;
         when "011010011111" => index <= 6;
         when "011010100000" => index <= 9;
         when "011010100001" => index <= 7;
         when "011010100010" => index <= 7;
         when "011010100011" => index <= 6;
         when "011010100100" => index <= 8;
         when "011010100101" => index <= 6;
         when "011010100110" => index <= 7;
         when "011010100111" => index <= 6;
         when "011010101000" => index <= 8;
         when "011010101001" => index <= 7;
         when "011010101010" => index <= 7;
         when "011010101011" => index <= 6;
         when "011010101100" => index <= 7;
         when "011010101101" => index <= 6;
         when "011010101110" => index <= 6;
         when "011010101111" => index <= 6;
         when "011010110000" => index <= 8;
         when "011010110001" => index <= 7;
         when "011010110010" => index <= 7;
         when "011010110011" => index <= 6;
         when "011010110100" => index <= 7;
         when "011010110101" => index <= 6;
         when "011010110110" => index <= 6;
         when "011010110111" => index <= 6;
         when "011010111000" => index <= 7;
         when "011010111001" => index <= 6;
         when "011010111010" => index <= 7;
         when "011010111011" => index <= 6;
         when "011010111100" => index <= 7;
         when "011010111101" => index <= 6;
         when "011010111110" => index <= 6;
         when "011010111111" => index <= 6;
         when "011011000000" => index <= 9;
         when "011011000001" => index <= 7;
         when "011011000010" => index <= 8;
         when "011011000011" => index <= 6;
         when "011011000100" => index <= 8;
         when "011011000101" => index <= 7;
         when "011011000110" => index <= 7;
         when "011011000111" => index <= 6;
         when "011011001000" => index <= 8;
         when "011011001001" => index <= 7;
         when "011011001010" => index <= 7;
         when "011011001011" => index <= 6;
         when "011011001100" => index <= 7;
         when "011011001101" => index <= 6;
         when "011011001110" => index <= 6;
         when "011011001111" => index <= 6;
         when "011011010000" => index <= 8;
         when "011011010001" => index <= 7;
         when "011011010010" => index <= 7;
         when "011011010011" => index <= 6;
         when "011011010100" => index <= 7;
         when "011011010101" => index <= 6;
         when "011011010110" => index <= 7;
         when "011011010111" => index <= 6;
         when "011011011000" => index <= 8;
         when "011011011001" => index <= 7;
         when "011011011010" => index <= 7;
         when "011011011011" => index <= 6;
         when "011011011100" => index <= 7;
         when "011011011101" => index <= 6;
         when "011011011110" => index <= 6;
         when "011011011111" => index <= 6;
         when "011011100000" => index <= 8;
         when "011011100001" => index <= 7;
         when "011011100010" => index <= 7;
         when "011011100011" => index <= 6;
         when "011011100100" => index <= 8;
         when "011011100101" => index <= 7;
         when "011011100110" => index <= 7;
         when "011011100111" => index <= 6;
         when "011011101000" => index <= 8;
         when "011011101001" => index <= 7;
         when "011011101010" => index <= 7;
         when "011011101011" => index <= 6;
         when "011011101100" => index <= 7;
         when "011011101101" => index <= 6;
         when "011011101110" => index <= 6;
         when "011011101111" => index <= 6;
         when "011011110000" => index <= 8;
         when "011011110001" => index <= 7;
         when "011011110010" => index <= 7;
         when "011011110011" => index <= 6;
         when "011011110100" => index <= 7;
         when "011011110101" => index <= 6;
         when "011011110110" => index <= 6;
         when "011011110111" => index <= 6;
         when "011011111000" => index <= 7;
         when "011011111001" => index <= 6;
         when "011011111010" => index <= 7;
         when "011011111011" => index <= 6;
         when "011011111100" => index <= 7;
         when "011011111101" => index <= 6;
         when "011011111110" => index <= 6;
         when "011011111111" => index <= 6;
         when "011100000000" => index <= 10;
         when "011100000001" => index <= 8;
         when "011100000010" => index <= 8;
         when "011100000011" => index <= 7;
         when "011100000100" => index <= 8;
         when "011100000101" => index <= 7;
         when "011100000110" => index <= 7;
         when "011100000111" => index <= 6;
         when "011100001000" => index <= 8;
         when "011100001001" => index <= 7;
         when "011100001010" => index <= 7;
         when "011100001011" => index <= 6;
         when "011100001100" => index <= 7;
         when "011100001101" => index <= 6;
         when "011100001110" => index <= 6;
         when "011100001111" => index <= 6;
         when "011100010000" => index <= 9;
         when "011100010001" => index <= 7;
         when "011100010010" => index <= 7;
         when "011100010011" => index <= 6;
         when "011100010100" => index <= 8;
         when "011100010101" => index <= 6;
         when "011100010110" => index <= 7;
         when "011100010111" => index <= 6;
         when "011100011000" => index <= 8;
         when "011100011001" => index <= 7;
         when "011100011010" => index <= 7;
         when "011100011011" => index <= 6;
         when "011100011100" => index <= 7;
         when "011100011101" => index <= 6;
         when "011100011110" => index <= 6;
         when "011100011111" => index <= 6;
         when "011100100000" => index <= 9;
         when "011100100001" => index <= 7;
         when "011100100010" => index <= 8;
         when "011100100011" => index <= 6;
         when "011100100100" => index <= 8;
         when "011100100101" => index <= 7;
         when "011100100110" => index <= 7;
         when "011100100111" => index <= 6;
         when "011100101000" => index <= 8;
         when "011100101001" => index <= 7;
         when "011100101010" => index <= 7;
         when "011100101011" => index <= 6;
         when "011100101100" => index <= 7;
         when "011100101101" => index <= 6;
         when "011100101110" => index <= 6;
         when "011100101111" => index <= 6;
         when "011100110000" => index <= 8;
         when "011100110001" => index <= 7;
         when "011100110010" => index <= 7;
         when "011100110011" => index <= 6;
         when "011100110100" => index <= 7;
         when "011100110101" => index <= 6;
         when "011100110110" => index <= 7;
         when "011100110111" => index <= 6;
         when "011100111000" => index <= 8;
         when "011100111001" => index <= 7;
         when "011100111010" => index <= 7;
         when "011100111011" => index <= 6;
         when "011100111100" => index <= 7;
         when "011100111101" => index <= 6;
         when "011100111110" => index <= 6;
         when "011100111111" => index <= 6;
         when "011101000000" => index <= 9;
         when "011101000001" => index <= 8;
         when "011101000010" => index <= 8;
         when "011101000011" => index <= 7;
         when "011101000100" => index <= 8;
         when "011101000101" => index <= 7;
         when "011101000110" => index <= 7;
         when "011101000111" => index <= 6;
         when "011101001000" => index <= 8;
         when "011101001001" => index <= 7;
         when "011101001010" => index <= 7;
         when "011101001011" => index <= 6;
         when "011101001100" => index <= 7;
         when "011101001101" => index <= 6;
         when "011101001110" => index <= 7;
         when "011101001111" => index <= 6;
         when "011101010000" => index <= 8;
         when "011101010001" => index <= 7;
         when "011101010010" => index <= 7;
         when "011101010011" => index <= 6;
         when "011101010100" => index <= 8;
         when "011101010101" => index <= 7;
         when "011101010110" => index <= 7;
         when "011101010111" => index <= 6;
         when "011101011000" => index <= 8;
         when "011101011001" => index <= 7;
         when "011101011010" => index <= 7;
         when "011101011011" => index <= 6;
         when "011101011100" => index <= 7;
         when "011101011101" => index <= 6;
         when "011101011110" => index <= 6;
         when "011101011111" => index <= 6;
         when "011101100000" => index <= 9;
         when "011101100001" => index <= 7;
         when "011101100010" => index <= 8;
         when "011101100011" => index <= 7;
         when "011101100100" => index <= 8;
         when "011101100101" => index <= 7;
         when "011101100110" => index <= 7;
         when "011101100111" => index <= 6;
         when "011101101000" => index <= 8;
         when "011101101001" => index <= 7;
         when "011101101010" => index <= 7;
         when "011101101011" => index <= 6;
         when "011101101100" => index <= 7;
         when "011101101101" => index <= 6;
         when "011101101110" => index <= 6;
         when "011101101111" => index <= 6;
         when "011101110000" => index <= 8;
         when "011101110001" => index <= 7;
         when "011101110010" => index <= 7;
         when "011101110011" => index <= 6;
         when "011101110100" => index <= 7;
         when "011101110101" => index <= 6;
         when "011101110110" => index <= 7;
         when "011101110111" => index <= 6;
         when "011101111000" => index <= 7;
         when "011101111001" => index <= 7;
         when "011101111010" => index <= 7;
         when "011101111011" => index <= 6;
         when "011101111100" => index <= 7;
         when "011101111101" => index <= 6;
         when "011101111110" => index <= 6;
         when "011101111111" => index <= 6;
         when "011110000000" => index <= 10;
         when "011110000001" => index <= 8;
         when "011110000010" => index <= 8;
         when "011110000011" => index <= 7;
         when "011110000100" => index <= 8;
         when "011110000101" => index <= 7;
         when "011110000110" => index <= 7;
         when "011110000111" => index <= 6;
         when "011110001000" => index <= 8;
         when "011110001001" => index <= 7;
         when "011110001010" => index <= 7;
         when "011110001011" => index <= 6;
         when "011110001100" => index <= 8;
         when "011110001101" => index <= 7;
         when "011110001110" => index <= 7;
         when "011110001111" => index <= 6;
         when "011110010000" => index <= 9;
         when "011110010001" => index <= 7;
         when "011110010010" => index <= 8;
         when "011110010011" => index <= 7;
         when "011110010100" => index <= 8;
         when "011110010101" => index <= 7;
         when "011110010110" => index <= 7;
         when "011110010111" => index <= 6;
         when "011110011000" => index <= 8;
         when "011110011001" => index <= 7;
         when "011110011010" => index <= 7;
         when "011110011011" => index <= 6;
         when "011110011100" => index <= 7;
         when "011110011101" => index <= 6;
         when "011110011110" => index <= 6;
         when "011110011111" => index <= 6;
         when "011110100000" => index <= 9;
         when "011110100001" => index <= 8;
         when "011110100010" => index <= 8;
         when "011110100011" => index <= 7;
         when "011110100100" => index <= 8;
         when "011110100101" => index <= 7;
         when "011110100110" => index <= 7;
         when "011110100111" => index <= 6;
         when "011110101000" => index <= 8;
         when "011110101001" => index <= 7;
         when "011110101010" => index <= 7;
         when "011110101011" => index <= 6;
         when "011110101100" => index <= 7;
         when "011110101101" => index <= 6;
         when "011110101110" => index <= 7;
         when "011110101111" => index <= 6;
         when "011110110000" => index <= 8;
         when "011110110001" => index <= 7;
         when "011110110010" => index <= 7;
         when "011110110011" => index <= 6;
         when "011110110100" => index <= 7;
         when "011110110101" => index <= 7;
         when "011110110110" => index <= 7;
         when "011110110111" => index <= 6;
         when "011110111000" => index <= 8;
         when "011110111001" => index <= 7;
         when "011110111010" => index <= 7;
         when "011110111011" => index <= 6;
         when "011110111100" => index <= 7;
         when "011110111101" => index <= 6;
         when "011110111110" => index <= 6;
         when "011110111111" => index <= 6;
         when "011111000000" => index <= 9;
         when "011111000001" => index <= 8;
         when "011111000010" => index <= 8;
         when "011111000011" => index <= 7;
         when "011111000100" => index <= 8;
         when "011111000101" => index <= 7;
         when "011111000110" => index <= 7;
         when "011111000111" => index <= 6;
         when "011111001000" => index <= 8;
         when "011111001001" => index <= 7;
         when "011111001010" => index <= 7;
         when "011111001011" => index <= 6;
         when "011111001100" => index <= 7;
         when "011111001101" => index <= 7;
         when "011111001110" => index <= 7;
         when "011111001111" => index <= 6;
         when "011111010000" => index <= 8;
         when "011111010001" => index <= 7;
         when "011111010010" => index <= 7;
         when "011111010011" => index <= 7;
         when "011111010100" => index <= 8;
         when "011111010101" => index <= 7;
         when "011111010110" => index <= 7;
         when "011111010111" => index <= 6;
         when "011111011000" => index <= 8;
         when "011111011001" => index <= 7;
         when "011111011010" => index <= 7;
         when "011111011011" => index <= 6;
         when "011111011100" => index <= 7;
         when "011111011101" => index <= 6;
         when "011111011110" => index <= 7;
         when "011111011111" => index <= 6;
         when "011111100000" => index <= 8;
         when "011111100001" => index <= 7;
         when "011111100010" => index <= 8;
         when "011111100011" => index <= 7;
         when "011111100100" => index <= 8;
         when "011111100101" => index <= 7;
         when "011111100110" => index <= 7;
         when "011111100111" => index <= 6;
         when "011111101000" => index <= 8;
         when "011111101001" => index <= 7;
         when "011111101010" => index <= 7;
         when "011111101011" => index <= 6;
         when "011111101100" => index <= 7;
         when "011111101101" => index <= 7;
         when "011111101110" => index <= 7;
         when "011111101111" => index <= 6;
         when "011111110000" => index <= 8;
         when "011111110001" => index <= 7;
         when "011111110010" => index <= 7;
         when "011111110011" => index <= 7;
         when "011111110100" => index <= 7;
         when "011111110101" => index <= 7;
         when "011111110110" => index <= 7;
         when "011111110111" => index <= 6;
         when "011111111000" => index <= 8;
         when "011111111001" => index <= 7;
         when "011111111010" => index <= 7;
         when "011111111011" => index <= 6;
         when "011111111100" => index <= 7;
         when "011111111101" => index <= 6;
         when "011111111110" => index <= 6;
         when "011111111111" => index <= 6;
         when "100000000000" => index <= 12;
         when "100000000001" => index <= 6;
         when "100000000010" => index <= 7;
         when "100000000011" => index <= 5;
         when "100000000100" => index <= 8;
         when "100000000101" => index <= 5;
         when "100000000110" => index <= 6;
         when "100000000111" => index <= 4;
         when "100000001000" => index <= 8;
         when "100000001001" => index <= 6;
         when "100000001010" => index <= 6;
         when "100000001011" => index <= 5;
         when "100000001100" => index <= 6;
         when "100000001101" => index <= 5;
         when "100000001110" => index <= 5;
         when "100000001111" => index <= 4;
         when "100000010000" => index <= 8;
         when "100000010001" => index <= 6;
         when "100000010010" => index <= 6;
         when "100000010011" => index <= 5;
         when "100000010100" => index <= 7;
         when "100000010101" => index <= 5;
         when "100000010110" => index <= 6;
         when "100000010111" => index <= 5;
         when "100000011000" => index <= 7;
         when "100000011001" => index <= 6;
         when "100000011010" => index <= 6;
         when "100000011011" => index <= 5;
         when "100000011100" => index <= 6;
         when "100000011101" => index <= 5;
         when "100000011110" => index <= 5;
         when "100000011111" => index <= 4;
         when "100000100000" => index <= 9;
         when "100000100001" => index <= 6;
         when "100000100010" => index <= 7;
         when "100000100011" => index <= 5;
         when "100000100100" => index <= 7;
         when "100000100101" => index <= 6;
         when "100000100110" => index <= 6;
         when "100000100111" => index <= 5;
         when "100000101000" => index <= 7;
         when "100000101001" => index <= 6;
         when "100000101010" => index <= 6;
         when "100000101011" => index <= 5;
         when "100000101100" => index <= 6;
         when "100000101101" => index <= 5;
         when "100000101110" => index <= 5;
         when "100000101111" => index <= 5;
         when "100000110000" => index <= 8;
         when "100000110001" => index <= 6;
         when "100000110010" => index <= 6;
         when "100000110011" => index <= 5;
         when "100000110100" => index <= 6;
         when "100000110101" => index <= 5;
         when "100000110110" => index <= 6;
         when "100000110111" => index <= 5;
         when "100000111000" => index <= 7;
         when "100000111001" => index <= 6;
         when "100000111010" => index <= 6;
         when "100000111011" => index <= 5;
         when "100000111100" => index <= 6;
         when "100000111101" => index <= 5;
         when "100000111110" => index <= 5;
         when "100000111111" => index <= 5;
         when "100001000000" => index <= 10;
         when "100001000001" => index <= 7;
         when "100001000010" => index <= 7;
         when "100001000011" => index <= 6;
         when "100001000100" => index <= 7;
         when "100001000101" => index <= 6;
         when "100001000110" => index <= 6;
         when "100001000111" => index <= 5;
         when "100001001000" => index <= 8;
         when "100001001001" => index <= 6;
         when "100001001010" => index <= 6;
         when "100001001011" => index <= 5;
         when "100001001100" => index <= 6;
         when "100001001101" => index <= 5;
         when "100001001110" => index <= 6;
         when "100001001111" => index <= 5;
         when "100001010000" => index <= 8;
         when "100001010001" => index <= 6;
         when "100001010010" => index <= 6;
         when "100001010011" => index <= 5;
         when "100001010100" => index <= 7;
         when "100001010101" => index <= 6;
         when "100001010110" => index <= 6;
         when "100001010111" => index <= 5;
         when "100001011000" => index <= 7;
         when "100001011001" => index <= 6;
         when "100001011010" => index <= 6;
         when "100001011011" => index <= 5;
         when "100001011100" => index <= 6;
         when "100001011101" => index <= 5;
         when "100001011110" => index <= 6;
         when "100001011111" => index <= 5;
         when "100001100000" => index <= 8;
         when "100001100001" => index <= 6;
         when "100001100010" => index <= 7;
         when "100001100011" => index <= 6;
         when "100001100100" => index <= 7;
         when "100001100101" => index <= 6;
         when "100001100110" => index <= 6;
         when "100001100111" => index <= 5;
         when "100001101000" => index <= 7;
         when "100001101001" => index <= 6;
         when "100001101010" => index <= 6;
         when "100001101011" => index <= 5;
         when "100001101100" => index <= 6;
         when "100001101101" => index <= 6;
         when "100001101110" => index <= 6;
         when "100001101111" => index <= 5;
         when "100001110000" => index <= 8;
         when "100001110001" => index <= 6;
         when "100001110010" => index <= 6;
         when "100001110011" => index <= 6;
         when "100001110100" => index <= 7;
         when "100001110101" => index <= 6;
         when "100001110110" => index <= 6;
         when "100001110111" => index <= 5;
         when "100001111000" => index <= 7;
         when "100001111001" => index <= 6;
         when "100001111010" => index <= 6;
         when "100001111011" => index <= 5;
         when "100001111100" => index <= 6;
         when "100001111101" => index <= 5;
         when "100001111110" => index <= 6;
         when "100001111111" => index <= 5;
         when "100010000000" => index <= 10;
         when "100010000001" => index <= 7;
         when "100010000010" => index <= 7;
         when "100010000011" => index <= 6;
         when "100010000100" => index <= 8;
         when "100010000101" => index <= 6;
         when "100010000110" => index <= 6;
         when "100010000111" => index <= 5;
         when "100010001000" => index <= 8;
         when "100010001001" => index <= 6;
         when "100010001010" => index <= 6;
         when "100010001011" => index <= 5;
         when "100010001100" => index <= 7;
         when "100010001101" => index <= 6;
         when "100010001110" => index <= 6;
         when "100010001111" => index <= 5;
         when "100010010000" => index <= 8;
         when "100010010001" => index <= 6;
         when "100010010010" => index <= 7;
         when "100010010011" => index <= 6;
         when "100010010100" => index <= 7;
         when "100010010101" => index <= 6;
         when "100010010110" => index <= 6;
         when "100010010111" => index <= 5;
         when "100010011000" => index <= 7;
         when "100010011001" => index <= 6;
         when "100010011010" => index <= 6;
         when "100010011011" => index <= 5;
         when "100010011100" => index <= 6;
         when "100010011101" => index <= 6;
         when "100010011110" => index <= 6;
         when "100010011111" => index <= 5;
         when "100010100000" => index <= 9;
         when "100010100001" => index <= 7;
         when "100010100010" => index <= 7;
         when "100010100011" => index <= 6;
         when "100010100100" => index <= 7;
         when "100010100101" => index <= 6;
         when "100010100110" => index <= 6;
         when "100010100111" => index <= 5;
         when "100010101000" => index <= 8;
         when "100010101001" => index <= 6;
         when "100010101010" => index <= 6;
         when "100010101011" => index <= 6;
         when "100010101100" => index <= 7;
         when "100010101101" => index <= 6;
         when "100010101110" => index <= 6;
         when "100010101111" => index <= 5;
         when "100010110000" => index <= 8;
         when "100010110001" => index <= 6;
         when "100010110010" => index <= 7;
         when "100010110011" => index <= 6;
         when "100010110100" => index <= 7;
         when "100010110101" => index <= 6;
         when "100010110110" => index <= 6;
         when "100010110111" => index <= 5;
         when "100010111000" => index <= 7;
         when "100010111001" => index <= 6;
         when "100010111010" => index <= 6;
         when "100010111011" => index <= 5;
         when "100010111100" => index <= 6;
         when "100010111101" => index <= 6;
         when "100010111110" => index <= 6;
         when "100010111111" => index <= 5;
         when "100011000000" => index <= 9;
         when "100011000001" => index <= 7;
         when "100011000010" => index <= 7;
         when "100011000011" => index <= 6;
         when "100011000100" => index <= 8;
         when "100011000101" => index <= 6;
         when "100011000110" => index <= 6;
         when "100011000111" => index <= 6;
         when "100011001000" => index <= 8;
         when "100011001001" => index <= 6;
         when "100011001010" => index <= 7;
         when "100011001011" => index <= 6;
         when "100011001100" => index <= 7;
         when "100011001101" => index <= 6;
         when "100011001110" => index <= 6;
         when "100011001111" => index <= 5;
         when "100011010000" => index <= 8;
         when "100011010001" => index <= 7;
         when "100011010010" => index <= 7;
         when "100011010011" => index <= 6;
         when "100011010100" => index <= 7;
         when "100011010101" => index <= 6;
         when "100011010110" => index <= 6;
         when "100011010111" => index <= 5;
         when "100011011000" => index <= 7;
         when "100011011001" => index <= 6;
         when "100011011010" => index <= 6;
         when "100011011011" => index <= 6;
         when "100011011100" => index <= 6;
         when "100011011101" => index <= 6;
         when "100011011110" => index <= 6;
         when "100011011111" => index <= 5;
         when "100011100000" => index <= 8;
         when "100011100001" => index <= 7;
         when "100011100010" => index <= 7;
         when "100011100011" => index <= 6;
         when "100011100100" => index <= 7;
         when "100011100101" => index <= 6;
         when "100011100110" => index <= 6;
         when "100011100111" => index <= 6;
         when "100011101000" => index <= 7;
         when "100011101001" => index <= 6;
         when "100011101010" => index <= 6;
         when "100011101011" => index <= 6;
         when "100011101100" => index <= 7;
         when "100011101101" => index <= 6;
         when "100011101110" => index <= 6;
         when "100011101111" => index <= 5;
         when "100011110000" => index <= 8;
         when "100011110001" => index <= 6;
         when "100011110010" => index <= 7;
         when "100011110011" => index <= 6;
         when "100011110100" => index <= 7;
         when "100011110101" => index <= 6;
         when "100011110110" => index <= 6;
         when "100011110111" => index <= 6;
         when "100011111000" => index <= 7;
         when "100011111001" => index <= 6;
         when "100011111010" => index <= 6;
         when "100011111011" => index <= 6;
         when "100011111100" => index <= 6;
         when "100011111101" => index <= 6;
         when "100011111110" => index <= 6;
         when "100011111111" => index <= 5;
         when "100100000000" => index <= 10;
         when "100100000001" => index <= 7;
         when "100100000010" => index <= 8;
         when "100100000011" => index <= 6;
         when "100100000100" => index <= 8;
         when "100100000101" => index <= 6;
         when "100100000110" => index <= 6;
         when "100100000111" => index <= 5;
         when "100100001000" => index <= 8;
         when "100100001001" => index <= 6;
         when "100100001010" => index <= 7;
         when "100100001011" => index <= 6;
         when "100100001100" => index <= 7;
         when "100100001101" => index <= 6;
         when "100100001110" => index <= 6;
         when "100100001111" => index <= 5;
         when "100100010000" => index <= 9;
         when "100100010001" => index <= 7;
         when "100100010010" => index <= 7;
         when "100100010011" => index <= 6;
         when "100100010100" => index <= 7;
         when "100100010101" => index <= 6;
         when "100100010110" => index <= 6;
         when "100100010111" => index <= 5;
         when "100100011000" => index <= 8;
         when "100100011001" => index <= 6;
         when "100100011010" => index <= 6;
         when "100100011011" => index <= 6;
         when "100100011100" => index <= 7;
         when "100100011101" => index <= 6;
         when "100100011110" => index <= 6;
         when "100100011111" => index <= 5;
         when "100100100000" => index <= 9;
         when "100100100001" => index <= 7;
         when "100100100010" => index <= 7;
         when "100100100011" => index <= 6;
         when "100100100100" => index <= 8;
         when "100100100101" => index <= 6;
         when "100100100110" => index <= 6;
         when "100100100111" => index <= 6;
         when "100100101000" => index <= 8;
         when "100100101001" => index <= 6;
         when "100100101010" => index <= 7;
         when "100100101011" => index <= 6;
         when "100100101100" => index <= 7;
         when "100100101101" => index <= 6;
         when "100100101110" => index <= 6;
         when "100100101111" => index <= 5;
         when "100100110000" => index <= 8;
         when "100100110001" => index <= 7;
         when "100100110010" => index <= 7;
         when "100100110011" => index <= 6;
         when "100100110100" => index <= 7;
         when "100100110101" => index <= 6;
         when "100100110110" => index <= 6;
         when "100100110111" => index <= 5;
         when "100100111000" => index <= 7;
         when "100100111001" => index <= 6;
         when "100100111010" => index <= 6;
         when "100100111011" => index <= 6;
         when "100100111100" => index <= 6;
         when "100100111101" => index <= 6;
         when "100100111110" => index <= 6;
         when "100100111111" => index <= 5;
         when "100101000000" => index <= 9;
         when "100101000001" => index <= 7;
         when "100101000010" => index <= 8;
         when "100101000011" => index <= 6;
         when "100101000100" => index <= 8;
         when "100101000101" => index <= 6;
         when "100101000110" => index <= 7;
         when "100101000111" => index <= 6;
         when "100101001000" => index <= 8;
         when "100101001001" => index <= 7;
         when "100101001010" => index <= 7;
         when "100101001011" => index <= 6;
         when "100101001100" => index <= 7;
         when "100101001101" => index <= 6;
         when "100101001110" => index <= 6;
         when "100101001111" => index <= 5;
         when "100101010000" => index <= 8;
         when "100101010001" => index <= 7;
         when "100101010010" => index <= 7;
         when "100101010011" => index <= 6;
         when "100101010100" => index <= 7;
         when "100101010101" => index <= 6;
         when "100101010110" => index <= 6;
         when "100101010111" => index <= 6;
         when "100101011000" => index <= 7;
         when "100101011001" => index <= 6;
         when "100101011010" => index <= 6;
         when "100101011011" => index <= 6;
         when "100101011100" => index <= 7;
         when "100101011101" => index <= 6;
         when "100101011110" => index <= 6;
         when "100101011111" => index <= 5;
         when "100101100000" => index <= 8;
         when "100101100001" => index <= 7;
         when "100101100010" => index <= 7;
         when "100101100011" => index <= 6;
         when "100101100100" => index <= 7;
         when "100101100101" => index <= 6;
         when "100101100110" => index <= 6;
         when "100101100111" => index <= 6;
         when "100101101000" => index <= 8;
         when "100101101001" => index <= 6;
         when "100101101010" => index <= 7;
         when "100101101011" => index <= 6;
         when "100101101100" => index <= 7;
         when "100101101101" => index <= 6;
         when "100101101110" => index <= 6;
         when "100101101111" => index <= 6;
         when "100101110000" => index <= 8;
         when "100101110001" => index <= 7;
         when "100101110010" => index <= 7;
         when "100101110011" => index <= 6;
         when "100101110100" => index <= 7;
         when "100101110101" => index <= 6;
         when "100101110110" => index <= 6;
         when "100101110111" => index <= 6;
         when "100101111000" => index <= 7;
         when "100101111001" => index <= 6;
         when "100101111010" => index <= 6;
         when "100101111011" => index <= 6;
         when "100101111100" => index <= 7;
         when "100101111101" => index <= 6;
         when "100101111110" => index <= 6;
         when "100101111111" => index <= 5;
         when "100110000000" => index <= 10;
         when "100110000001" => index <= 8;
         when "100110000010" => index <= 8;
         when "100110000011" => index <= 6;
         when "100110000100" => index <= 8;
         when "100110000101" => index <= 7;
         when "100110000110" => index <= 7;
         when "100110000111" => index <= 6;
         when "100110001000" => index <= 8;
         when "100110001001" => index <= 7;
         when "100110001010" => index <= 7;
         when "100110001011" => index <= 6;
         when "100110001100" => index <= 7;
         when "100110001101" => index <= 6;
         when "100110001110" => index <= 6;
         when "100110001111" => index <= 6;
         when "100110010000" => index <= 8;
         when "100110010001" => index <= 7;
         when "100110010010" => index <= 7;
         when "100110010011" => index <= 6;
         when "100110010100" => index <= 7;
         when "100110010101" => index <= 6;
         when "100110010110" => index <= 6;
         when "100110010111" => index <= 6;
         when "100110011000" => index <= 8;
         when "100110011001" => index <= 6;
         when "100110011010" => index <= 7;
         when "100110011011" => index <= 6;
         when "100110011100" => index <= 7;
         when "100110011101" => index <= 6;
         when "100110011110" => index <= 6;
         when "100110011111" => index <= 6;
         when "100110100000" => index <= 9;
         when "100110100001" => index <= 7;
         when "100110100010" => index <= 7;
         when "100110100011" => index <= 6;
         when "100110100100" => index <= 8;
         when "100110100101" => index <= 6;
         when "100110100110" => index <= 7;
         when "100110100111" => index <= 6;
         when "100110101000" => index <= 8;
         when "100110101001" => index <= 7;
         when "100110101010" => index <= 7;
         when "100110101011" => index <= 6;
         when "100110101100" => index <= 7;
         when "100110101101" => index <= 6;
         when "100110101110" => index <= 6;
         when "100110101111" => index <= 6;
         when "100110110000" => index <= 8;
         when "100110110001" => index <= 7;
         when "100110110010" => index <= 7;
         when "100110110011" => index <= 6;
         when "100110110100" => index <= 7;
         when "100110110101" => index <= 6;
         when "100110110110" => index <= 6;
         when "100110110111" => index <= 6;
         when "100110111000" => index <= 7;
         when "100110111001" => index <= 6;
         when "100110111010" => index <= 7;
         when "100110111011" => index <= 6;
         when "100110111100" => index <= 7;
         when "100110111101" => index <= 6;
         when "100110111110" => index <= 6;
         when "100110111111" => index <= 6;
         when "100111000000" => index <= 9;
         when "100111000001" => index <= 7;
         when "100111000010" => index <= 8;
         when "100111000011" => index <= 6;
         when "100111000100" => index <= 8;
         when "100111000101" => index <= 7;
         when "100111000110" => index <= 7;
         when "100111000111" => index <= 6;
         when "100111001000" => index <= 8;
         when "100111001001" => index <= 7;
         when "100111001010" => index <= 7;
         when "100111001011" => index <= 6;
         when "100111001100" => index <= 7;
         when "100111001101" => index <= 6;
         when "100111001110" => index <= 6;
         when "100111001111" => index <= 6;
         when "100111010000" => index <= 8;
         when "100111010001" => index <= 7;
         when "100111010010" => index <= 7;
         when "100111010011" => index <= 6;
         when "100111010100" => index <= 7;
         when "100111010101" => index <= 6;
         when "100111010110" => index <= 7;
         when "100111010111" => index <= 6;
         when "100111011000" => index <= 8;
         when "100111011001" => index <= 7;
         when "100111011010" => index <= 7;
         when "100111011011" => index <= 6;
         when "100111011100" => index <= 7;
         when "100111011101" => index <= 6;
         when "100111011110" => index <= 6;
         when "100111011111" => index <= 6;
         when "100111100000" => index <= 8;
         when "100111100001" => index <= 7;
         when "100111100010" => index <= 7;
         when "100111100011" => index <= 6;
         when "100111100100" => index <= 8;
         when "100111100101" => index <= 7;
         when "100111100110" => index <= 7;
         when "100111100111" => index <= 6;
         when "100111101000" => index <= 8;
         when "100111101001" => index <= 7;
         when "100111101010" => index <= 7;
         when "100111101011" => index <= 6;
         when "100111101100" => index <= 7;
         when "100111101101" => index <= 6;
         when "100111101110" => index <= 6;
         when "100111101111" => index <= 6;
         when "100111110000" => index <= 8;
         when "100111110001" => index <= 7;
         when "100111110010" => index <= 7;
         when "100111110011" => index <= 6;
         when "100111110100" => index <= 7;
         when "100111110101" => index <= 6;
         when "100111110110" => index <= 6;
         when "100111110111" => index <= 6;
         when "100111111000" => index <= 7;
         when "100111111001" => index <= 6;
         when "100111111010" => index <= 7;
         when "100111111011" => index <= 6;
         when "100111111100" => index <= 7;
         when "100111111101" => index <= 6;
         when "100111111110" => index <= 6;
         when "100111111111" => index <= 6;
         when "101000000000" => index <= 11;
         when "101000000001" => index <= 8;
         when "101000000010" => index <= 8;
         when "101000000011" => index <= 6;
         when "101000000100" => index <= 8;
         when "101000000101" => index <= 6;
         when "101000000110" => index <= 7;
         when "101000000111" => index <= 6;
         when "101000001000" => index <= 9;
         when "101000001001" => index <= 7;
         when "101000001010" => index <= 7;
         when "101000001011" => index <= 6;
         when "101000001100" => index <= 7;
         when "101000001101" => index <= 6;
         when "101000001110" => index <= 6;
         when "101000001111" => index <= 5;
         when "101000010000" => index <= 9;
         when "101000010001" => index <= 7;
         when "101000010010" => index <= 7;
         when "101000010011" => index <= 6;
         when "101000010100" => index <= 8;
         when "101000010101" => index <= 6;
         when "101000010110" => index <= 6;
         when "101000010111" => index <= 6;
         when "101000011000" => index <= 8;
         when "101000011001" => index <= 6;
         when "101000011010" => index <= 7;
         when "101000011011" => index <= 6;
         when "101000011100" => index <= 7;
         when "101000011101" => index <= 6;
         when "101000011110" => index <= 6;
         when "101000011111" => index <= 5;
         when "101000100000" => index <= 9;
         when "101000100001" => index <= 7;
         when "101000100010" => index <= 8;
         when "101000100011" => index <= 6;
         when "101000100100" => index <= 8;
         when "101000100101" => index <= 6;
         when "101000100110" => index <= 7;
         when "101000100111" => index <= 6;
         when "101000101000" => index <= 8;
         when "101000101001" => index <= 7;
         when "101000101010" => index <= 7;
         when "101000101011" => index <= 6;
         when "101000101100" => index <= 7;
         when "101000101101" => index <= 6;
         when "101000101110" => index <= 6;
         when "101000101111" => index <= 5;
         when "101000110000" => index <= 8;
         when "101000110001" => index <= 7;
         when "101000110010" => index <= 7;
         when "101000110011" => index <= 6;
         when "101000110100" => index <= 7;
         when "101000110101" => index <= 6;
         when "101000110110" => index <= 6;
         when "101000110111" => index <= 6;
         when "101000111000" => index <= 7;
         when "101000111001" => index <= 6;
         when "101000111010" => index <= 6;
         when "101000111011" => index <= 6;
         when "101000111100" => index <= 7;
         when "101000111101" => index <= 6;
         when "101000111110" => index <= 6;
         when "101000111111" => index <= 5;
         when "101001000000" => index <= 10;
         when "101001000001" => index <= 8;
         when "101001000010" => index <= 8;
         when "101001000011" => index <= 6;
         when "101001000100" => index <= 8;
         when "101001000101" => index <= 7;
         when "101001000110" => index <= 7;
         when "101001000111" => index <= 6;
         when "101001001000" => index <= 8;
         when "101001001001" => index <= 7;
         when "101001001010" => index <= 7;
         when "101001001011" => index <= 6;
         when "101001001100" => index <= 7;
         when "101001001101" => index <= 6;
         when "101001001110" => index <= 6;
         when "101001001111" => index <= 6;
         when "101001010000" => index <= 8;
         when "101001010001" => index <= 7;
         when "101001010010" => index <= 7;
         when "101001010011" => index <= 6;
         when "101001010100" => index <= 7;
         when "101001010101" => index <= 6;
         when "101001010110" => index <= 6;
         when "101001010111" => index <= 6;
         when "101001011000" => index <= 8;
         when "101001011001" => index <= 6;
         when "101001011010" => index <= 7;
         when "101001011011" => index <= 6;
         when "101001011100" => index <= 7;
         when "101001011101" => index <= 6;
         when "101001011110" => index <= 6;
         when "101001011111" => index <= 6;
         when "101001100000" => index <= 9;
         when "101001100001" => index <= 7;
         when "101001100010" => index <= 7;
         when "101001100011" => index <= 6;
         when "101001100100" => index <= 8;
         when "101001100101" => index <= 6;
         when "101001100110" => index <= 7;
         when "101001100111" => index <= 6;
         when "101001101000" => index <= 8;
         when "101001101001" => index <= 7;
         when "101001101010" => index <= 7;
         when "101001101011" => index <= 6;
         when "101001101100" => index <= 7;
         when "101001101101" => index <= 6;
         when "101001101110" => index <= 6;
         when "101001101111" => index <= 6;
         when "101001110000" => index <= 8;
         when "101001110001" => index <= 7;
         when "101001110010" => index <= 7;
         when "101001110011" => index <= 6;
         when "101001110100" => index <= 7;
         when "101001110101" => index <= 6;
         when "101001110110" => index <= 6;
         when "101001110111" => index <= 6;
         when "101001111000" => index <= 7;
         when "101001111001" => index <= 6;
         when "101001111010" => index <= 7;
         when "101001111011" => index <= 6;
         when "101001111100" => index <= 7;
         when "101001111101" => index <= 6;
         when "101001111110" => index <= 6;
         when "101001111111" => index <= 6;
         when "101010000000" => index <= 10;
         when "101010000001" => index <= 8;
         when "101010000010" => index <= 8;
         when "101010000011" => index <= 7;
         when "101010000100" => index <= 8;
         when "101010000101" => index <= 7;
         when "101010000110" => index <= 7;
         when "101010000111" => index <= 6;
         when "101010001000" => index <= 8;
         when "101010001001" => index <= 7;
         when "101010001010" => index <= 7;
         when "101010001011" => index <= 6;
         when "101010001100" => index <= 7;
         when "101010001101" => index <= 6;
         when "101010001110" => index <= 6;
         when "101010001111" => index <= 6;
         when "101010010000" => index <= 9;
         when "101010010001" => index <= 7;
         when "101010010010" => index <= 7;
         when "101010010011" => index <= 6;
         when "101010010100" => index <= 8;
         when "101010010101" => index <= 6;
         when "101010010110" => index <= 7;
         when "101010010111" => index <= 6;
         when "101010011000" => index <= 8;
         when "101010011001" => index <= 7;
         when "101010011010" => index <= 7;
         when "101010011011" => index <= 6;
         when "101010011100" => index <= 7;
         when "101010011101" => index <= 6;
         when "101010011110" => index <= 6;
         when "101010011111" => index <= 6;
         when "101010100000" => index <= 9;
         when "101010100001" => index <= 7;
         when "101010100010" => index <= 8;
         when "101010100011" => index <= 6;
         when "101010100100" => index <= 8;
         when "101010100101" => index <= 7;
         when "101010100110" => index <= 7;
         when "101010100111" => index <= 6;
         when "101010101000" => index <= 8;
         when "101010101001" => index <= 7;
         when "101010101010" => index <= 7;
         when "101010101011" => index <= 6;
         when "101010101100" => index <= 7;
         when "101010101101" => index <= 6;
         when "101010101110" => index <= 6;
         when "101010101111" => index <= 6;
         when "101010110000" => index <= 8;
         when "101010110001" => index <= 7;
         when "101010110010" => index <= 7;
         when "101010110011" => index <= 6;
         when "101010110100" => index <= 7;
         when "101010110101" => index <= 6;
         when "101010110110" => index <= 7;
         when "101010110111" => index <= 6;
         when "101010111000" => index <= 8;
         when "101010111001" => index <= 7;
         when "101010111010" => index <= 7;
         when "101010111011" => index <= 6;
         when "101010111100" => index <= 7;
         when "101010111101" => index <= 6;
         when "101010111110" => index <= 6;
         when "101010111111" => index <= 6;
         when "101011000000" => index <= 9;
         when "101011000001" => index <= 8;
         when "101011000010" => index <= 8;
         when "101011000011" => index <= 7;
         when "101011000100" => index <= 8;
         when "101011000101" => index <= 7;
         when "101011000110" => index <= 7;
         when "101011000111" => index <= 6;
         when "101011001000" => index <= 8;
         when "101011001001" => index <= 7;
         when "101011001010" => index <= 7;
         when "101011001011" => index <= 6;
         when "101011001100" => index <= 7;
         when "101011001101" => index <= 6;
         when "101011001110" => index <= 7;
         when "101011001111" => index <= 6;
         when "101011010000" => index <= 8;
         when "101011010001" => index <= 7;
         when "101011010010" => index <= 7;
         when "101011010011" => index <= 6;
         when "101011010100" => index <= 8;
         when "101011010101" => index <= 7;
         when "101011010110" => index <= 7;
         when "101011010111" => index <= 6;
         when "101011011000" => index <= 8;
         when "101011011001" => index <= 7;
         when "101011011010" => index <= 7;
         when "101011011011" => index <= 6;
         when "101011011100" => index <= 7;
         when "101011011101" => index <= 6;
         when "101011011110" => index <= 6;
         when "101011011111" => index <= 6;
         when "101011100000" => index <= 9;
         when "101011100001" => index <= 7;
         when "101011100010" => index <= 8;
         when "101011100011" => index <= 7;
         when "101011100100" => index <= 8;
         when "101011100101" => index <= 7;
         when "101011100110" => index <= 7;
         when "101011100111" => index <= 6;
         when "101011101000" => index <= 8;
         when "101011101001" => index <= 7;
         when "101011101010" => index <= 7;
         when "101011101011" => index <= 6;
         when "101011101100" => index <= 7;
         when "101011101101" => index <= 6;
         when "101011101110" => index <= 6;
         when "101011101111" => index <= 6;
         when "101011110000" => index <= 8;
         when "101011110001" => index <= 7;
         when "101011110010" => index <= 7;
         when "101011110011" => index <= 6;
         when "101011110100" => index <= 7;
         when "101011110101" => index <= 6;
         when "101011110110" => index <= 7;
         when "101011110111" => index <= 6;
         when "101011111000" => index <= 7;
         when "101011111001" => index <= 7;
         when "101011111010" => index <= 7;
         when "101011111011" => index <= 6;
         when "101011111100" => index <= 7;
         when "101011111101" => index <= 6;
         when "101011111110" => index <= 6;
         when "101011111111" => index <= 6;
         when "101100000000" => index <= 10;
         when "101100000001" => index <= 8;
         when "101100000010" => index <= 8;
         when "101100000011" => index <= 7;
         when "101100000100" => index <= 8;
         when "101100000101" => index <= 7;
         when "101100000110" => index <= 7;
         when "101100000111" => index <= 6;
         when "101100001000" => index <= 9;
         when "101100001001" => index <= 7;
         when "101100001010" => index <= 7;
         when "101100001011" => index <= 6;
         when "101100001100" => index <= 8;
         when "101100001101" => index <= 6;
         when "101100001110" => index <= 7;
         when "101100001111" => index <= 6;
         when "101100010000" => index <= 9;
         when "101100010001" => index <= 7;
         when "101100010010" => index <= 8;
         when "101100010011" => index <= 6;
         when "101100010100" => index <= 8;
         when "101100010101" => index <= 7;
         when "101100010110" => index <= 7;
         when "101100010111" => index <= 6;
         when "101100011000" => index <= 8;
         when "101100011001" => index <= 7;
         when "101100011010" => index <= 7;
         when "101100011011" => index <= 6;
         when "101100011100" => index <= 7;
         when "101100011101" => index <= 6;
         when "101100011110" => index <= 6;
         when "101100011111" => index <= 6;
         when "101100100000" => index <= 9;
         when "101100100001" => index <= 8;
         when "101100100010" => index <= 8;
         when "101100100011" => index <= 7;
         when "101100100100" => index <= 8;
         when "101100100101" => index <= 7;
         when "101100100110" => index <= 7;
         when "101100100111" => index <= 6;
         when "101100101000" => index <= 8;
         when "101100101001" => index <= 7;
         when "101100101010" => index <= 7;
         when "101100101011" => index <= 6;
         when "101100101100" => index <= 7;
         when "101100101101" => index <= 6;
         when "101100101110" => index <= 7;
         when "101100101111" => index <= 6;
         when "101100110000" => index <= 8;
         when "101100110001" => index <= 7;
         when "101100110010" => index <= 7;
         when "101100110011" => index <= 6;
         when "101100110100" => index <= 8;
         when "101100110101" => index <= 7;
         when "101100110110" => index <= 7;
         when "101100110111" => index <= 6;
         when "101100111000" => index <= 8;
         when "101100111001" => index <= 7;
         when "101100111010" => index <= 7;
         when "101100111011" => index <= 6;
         when "101100111100" => index <= 7;
         when "101100111101" => index <= 6;
         when "101100111110" => index <= 6;
         when "101100111111" => index <= 6;
         when "101101000000" => index <= 10;
         when "101101000001" => index <= 8;
         when "101101000010" => index <= 8;
         when "101101000011" => index <= 7;
         when "101101000100" => index <= 8;
         when "101101000101" => index <= 7;
         when "101101000110" => index <= 7;
         when "101101000111" => index <= 6;
         when "101101001000" => index <= 8;
         when "101101001001" => index <= 7;
         when "101101001010" => index <= 7;
         when "101101001011" => index <= 6;
         when "101101001100" => index <= 8;
         when "101101001101" => index <= 7;
         when "101101001110" => index <= 7;
         when "101101001111" => index <= 6;
         when "101101010000" => index <= 9;
         when "101101010001" => index <= 7;
         when "101101010010" => index <= 8;
         when "101101010011" => index <= 7;
         when "101101010100" => index <= 8;
         when "101101010101" => index <= 7;
         when "101101010110" => index <= 7;
         when "101101010111" => index <= 6;
         when "101101011000" => index <= 8;
         when "101101011001" => index <= 7;
         when "101101011010" => index <= 7;
         when "101101011011" => index <= 6;
         when "101101011100" => index <= 7;
         when "101101011101" => index <= 6;
         when "101101011110" => index <= 6;
         when "101101011111" => index <= 6;
         when "101101100000" => index <= 9;
         when "101101100001" => index <= 8;
         when "101101100010" => index <= 8;
         when "101101100011" => index <= 7;
         when "101101100100" => index <= 8;
         when "101101100101" => index <= 7;
         when "101101100110" => index <= 7;
         when "101101100111" => index <= 6;
         when "101101101000" => index <= 8;
         when "101101101001" => index <= 7;
         when "101101101010" => index <= 7;
         when "101101101011" => index <= 6;
         when "101101101100" => index <= 7;
         when "101101101101" => index <= 6;
         when "101101101110" => index <= 7;
         when "101101101111" => index <= 6;
         when "101101110000" => index <= 8;
         when "101101110001" => index <= 7;
         when "101101110010" => index <= 7;
         when "101101110011" => index <= 6;
         when "101101110100" => index <= 7;
         when "101101110101" => index <= 7;
         when "101101110110" => index <= 7;
         when "101101110111" => index <= 6;
         when "101101111000" => index <= 8;
         when "101101111001" => index <= 7;
         when "101101111010" => index <= 7;
         when "101101111011" => index <= 6;
         when "101101111100" => index <= 7;
         when "101101111101" => index <= 6;
         when "101101111110" => index <= 6;
         when "101101111111" => index <= 6;
         when "101110000000" => index <= 10;
         when "101110000001" => index <= 8;
         when "101110000010" => index <= 8;
         when "101110000011" => index <= 7;
         when "101110000100" => index <= 8;
         when "101110000101" => index <= 7;
         when "101110000110" => index <= 7;
         when "101110000111" => index <= 6;
         when "101110001000" => index <= 9;
         when "101110001001" => index <= 7;
         when "101110001010" => index <= 8;
         when "101110001011" => index <= 7;
         when "101110001100" => index <= 8;
         when "101110001101" => index <= 7;
         when "101110001110" => index <= 7;
         when "101110001111" => index <= 6;
         when "101110010000" => index <= 9;
         when "101110010001" => index <= 8;
         when "101110010010" => index <= 8;
         when "101110010011" => index <= 7;
         when "101110010100" => index <= 8;
         when "101110010101" => index <= 7;
         when "101110010110" => index <= 7;
         when "101110010111" => index <= 6;
         when "101110011000" => index <= 8;
         when "101110011001" => index <= 7;
         when "101110011010" => index <= 7;
         when "101110011011" => index <= 6;
         when "101110011100" => index <= 7;
         when "101110011101" => index <= 6;
         when "101110011110" => index <= 7;
         when "101110011111" => index <= 6;
         when "101110100000" => index <= 9;
         when "101110100001" => index <= 8;
         when "101110100010" => index <= 8;
         when "101110100011" => index <= 7;
         when "101110100100" => index <= 8;
         when "101110100101" => index <= 7;
         when "101110100110" => index <= 7;
         when "101110100111" => index <= 6;
         when "101110101000" => index <= 8;
         when "101110101001" => index <= 7;
         when "101110101010" => index <= 7;
         when "101110101011" => index <= 6;
         when "101110101100" => index <= 7;
         when "101110101101" => index <= 7;
         when "101110101110" => index <= 7;
         when "101110101111" => index <= 6;
         when "101110110000" => index <= 8;
         when "101110110001" => index <= 7;
         when "101110110010" => index <= 7;
         when "101110110011" => index <= 7;
         when "101110110100" => index <= 8;
         when "101110110101" => index <= 7;
         when "101110110110" => index <= 7;
         when "101110110111" => index <= 6;
         when "101110111000" => index <= 8;
         when "101110111001" => index <= 7;
         when "101110111010" => index <= 7;
         when "101110111011" => index <= 6;
         when "101110111100" => index <= 7;
         when "101110111101" => index <= 6;
         when "101110111110" => index <= 7;
         when "101110111111" => index <= 6;
         when "101111000000" => index <= 9;
         when "101111000001" => index <= 8;
         when "101111000010" => index <= 8;
         when "101111000011" => index <= 7;
         when "101111000100" => index <= 8;
         when "101111000101" => index <= 7;
         when "101111000110" => index <= 7;
         when "101111000111" => index <= 6;
         when "101111001000" => index <= 8;
         when "101111001001" => index <= 7;
         when "101111001010" => index <= 7;
         when "101111001011" => index <= 7;
         when "101111001100" => index <= 8;
         when "101111001101" => index <= 7;
         when "101111001110" => index <= 7;
         when "101111001111" => index <= 6;
         when "101111010000" => index <= 8;
         when "101111010001" => index <= 7;
         when "101111010010" => index <= 8;
         when "101111010011" => index <= 7;
         when "101111010100" => index <= 8;
         when "101111010101" => index <= 7;
         when "101111010110" => index <= 7;
         when "101111010111" => index <= 6;
         when "101111011000" => index <= 8;
         when "101111011001" => index <= 7;
         when "101111011010" => index <= 7;
         when "101111011011" => index <= 6;
         when "101111011100" => index <= 7;
         when "101111011101" => index <= 7;
         when "101111011110" => index <= 7;
         when "101111011111" => index <= 6;
         when "101111100000" => index <= 9;
         when "101111100001" => index <= 8;
         when "101111100010" => index <= 8;
         when "101111100011" => index <= 7;
         when "101111100100" => index <= 8;
         when "101111100101" => index <= 7;
         when "101111100110" => index <= 7;
         when "101111100111" => index <= 6;
         when "101111101000" => index <= 8;
         when "101111101001" => index <= 7;
         when "101111101010" => index <= 7;
         when "101111101011" => index <= 7;
         when "101111101100" => index <= 7;
         when "101111101101" => index <= 7;
         when "101111101110" => index <= 7;
         when "101111101111" => index <= 6;
         when "101111110000" => index <= 8;
         when "101111110001" => index <= 7;
         when "101111110010" => index <= 7;
         when "101111110011" => index <= 7;
         when "101111110100" => index <= 8;
         when "101111110101" => index <= 7;
         when "101111110110" => index <= 7;
         when "101111110111" => index <= 6;
         when "101111111000" => index <= 8;
         when "101111111001" => index <= 7;
         when "101111111010" => index <= 7;
         when "101111111011" => index <= 6;
         when "101111111100" => index <= 7;
         when "101111111101" => index <= 6;
         when "101111111110" => index <= 7;
         when "101111111111" => index <= 6;
         when "110000000000" => index <= 12;
         when "110000000001" => index <= 8;
         when "110000000010" => index <= 8;
         when "110000000011" => index <= 6;
         when "110000000100" => index <= 9;
         when "110000000101" => index <= 7;
         when "110000000110" => index <= 7;
         when "110000000111" => index <= 6;
         when "110000001000" => index <= 9;
         when "110000001001" => index <= 7;
         when "110000001010" => index <= 7;
         when "110000001011" => index <= 6;
         when "110000001100" => index <= 8;
         when "110000001101" => index <= 6;
         when "110000001110" => index <= 6;
         when "110000001111" => index <= 6;
         when "110000010000" => index <= 9;
         when "110000010001" => index <= 7;
         when "110000010010" => index <= 8;
         when "110000010011" => index <= 6;
         when "110000010100" => index <= 8;
         when "110000010101" => index <= 6;
         when "110000010110" => index <= 7;
         when "110000010111" => index <= 6;
         when "110000011000" => index <= 8;
         when "110000011001" => index <= 7;
         when "110000011010" => index <= 7;
         when "110000011011" => index <= 6;
         when "110000011100" => index <= 7;
         when "110000011101" => index <= 6;
         when "110000011110" => index <= 6;
         when "110000011111" => index <= 5;
         when "110000100000" => index <= 10;
         when "110000100001" => index <= 8;
         when "110000100010" => index <= 8;
         when "110000100011" => index <= 6;
         when "110000100100" => index <= 8;
         when "110000100101" => index <= 7;
         when "110000100110" => index <= 7;
         when "110000100111" => index <= 6;
         when "110000101000" => index <= 8;
         when "110000101001" => index <= 7;
         when "110000101010" => index <= 7;
         when "110000101011" => index <= 6;
         when "110000101100" => index <= 7;
         when "110000101101" => index <= 6;
         when "110000101110" => index <= 6;
         when "110000101111" => index <= 6;
         when "110000110000" => index <= 8;
         when "110000110001" => index <= 7;
         when "110000110010" => index <= 7;
         when "110000110011" => index <= 6;
         when "110000110100" => index <= 7;
         when "110000110101" => index <= 6;
         when "110000110110" => index <= 6;
         when "110000110111" => index <= 6;
         when "110000111000" => index <= 8;
         when "110000111001" => index <= 6;
         when "110000111010" => index <= 7;
         when "110000111011" => index <= 6;
         when "110000111100" => index <= 7;
         when "110000111101" => index <= 6;
         when "110000111110" => index <= 6;
         when "110000111111" => index <= 6;
         when "110001000000" => index <= 10;
         when "110001000001" => index <= 8;
         when "110001000010" => index <= 8;
         when "110001000011" => index <= 7;
         when "110001000100" => index <= 8;
         when "110001000101" => index <= 7;
         when "110001000110" => index <= 7;
         when "110001000111" => index <= 6;
         when "110001001000" => index <= 8;
         when "110001001001" => index <= 7;
         when "110001001010" => index <= 7;
         when "110001001011" => index <= 6;
         when "110001001100" => index <= 7;
         when "110001001101" => index <= 6;
         when "110001001110" => index <= 6;
         when "110001001111" => index <= 6;
         when "110001010000" => index <= 9;
         when "110001010001" => index <= 7;
         when "110001010010" => index <= 7;
         when "110001010011" => index <= 6;
         when "110001010100" => index <= 8;
         when "110001010101" => index <= 6;
         when "110001010110" => index <= 7;
         when "110001010111" => index <= 6;
         when "110001011000" => index <= 8;
         when "110001011001" => index <= 7;
         when "110001011010" => index <= 7;
         when "110001011011" => index <= 6;
         when "110001011100" => index <= 7;
         when "110001011101" => index <= 6;
         when "110001011110" => index <= 6;
         when "110001011111" => index <= 6;
         when "110001100000" => index <= 9;
         when "110001100001" => index <= 7;
         when "110001100010" => index <= 8;
         when "110001100011" => index <= 6;
         when "110001100100" => index <= 8;
         when "110001100101" => index <= 7;
         when "110001100110" => index <= 7;
         when "110001100111" => index <= 6;
         when "110001101000" => index <= 8;
         when "110001101001" => index <= 7;
         when "110001101010" => index <= 7;
         when "110001101011" => index <= 6;
         when "110001101100" => index <= 7;
         when "110001101101" => index <= 6;
         when "110001101110" => index <= 6;
         when "110001101111" => index <= 6;
         when "110001110000" => index <= 8;
         when "110001110001" => index <= 7;
         when "110001110010" => index <= 7;
         when "110001110011" => index <= 6;
         when "110001110100" => index <= 7;
         when "110001110101" => index <= 6;
         when "110001110110" => index <= 7;
         when "110001110111" => index <= 6;
         when "110001111000" => index <= 8;
         when "110001111001" => index <= 7;
         when "110001111010" => index <= 7;
         when "110001111011" => index <= 6;
         when "110001111100" => index <= 7;
         when "110001111101" => index <= 6;
         when "110001111110" => index <= 6;
         when "110001111111" => index <= 6;
         when "110010000000" => index <= 10;
         when "110010000001" => index <= 8;
         when "110010000010" => index <= 8;
         when "110010000011" => index <= 7;
         when "110010000100" => index <= 8;
         when "110010000101" => index <= 7;
         when "110010000110" => index <= 7;
         when "110010000111" => index <= 6;
         when "110010001000" => index <= 9;
         when "110010001001" => index <= 7;
         when "110010001010" => index <= 7;
         when "110010001011" => index <= 6;
         when "110010001100" => index <= 8;
         when "110010001101" => index <= 6;
         when "110010001110" => index <= 7;
         when "110010001111" => index <= 6;
         when "110010010000" => index <= 9;
         when "110010010001" => index <= 7;
         when "110010010010" => index <= 8;
         when "110010010011" => index <= 6;
         when "110010010100" => index <= 8;
         when "110010010101" => index <= 7;
         when "110010010110" => index <= 7;
         when "110010010111" => index <= 6;
         when "110010011000" => index <= 8;
         when "110010011001" => index <= 7;
         when "110010011010" => index <= 7;
         when "110010011011" => index <= 6;
         when "110010011100" => index <= 7;
         when "110010011101" => index <= 6;
         when "110010011110" => index <= 6;
         when "110010011111" => index <= 6;
         when "110010100000" => index <= 9;
         when "110010100001" => index <= 8;
         when "110010100010" => index <= 8;
         when "110010100011" => index <= 7;
         when "110010100100" => index <= 8;
         when "110010100101" => index <= 7;
         when "110010100110" => index <= 7;
         when "110010100111" => index <= 6;
         when "110010101000" => index <= 8;
         when "110010101001" => index <= 7;
         when "110010101010" => index <= 7;
         when "110010101011" => index <= 6;
         when "110010101100" => index <= 7;
         when "110010101101" => index <= 6;
         when "110010101110" => index <= 7;
         when "110010101111" => index <= 6;
         when "110010110000" => index <= 8;
         when "110010110001" => index <= 7;
         when "110010110010" => index <= 7;
         when "110010110011" => index <= 6;
         when "110010110100" => index <= 8;
         when "110010110101" => index <= 7;
         when "110010110110" => index <= 7;
         when "110010110111" => index <= 6;
         when "110010111000" => index <= 8;
         when "110010111001" => index <= 7;
         when "110010111010" => index <= 7;
         when "110010111011" => index <= 6;
         when "110010111100" => index <= 7;
         when "110010111101" => index <= 6;
         when "110010111110" => index <= 6;
         when "110010111111" => index <= 6;
         when "110011000000" => index <= 10;
         when "110011000001" => index <= 8;
         when "110011000010" => index <= 8;
         when "110011000011" => index <= 7;
         when "110011000100" => index <= 8;
         when "110011000101" => index <= 7;
         when "110011000110" => index <= 7;
         when "110011000111" => index <= 6;
         when "110011001000" => index <= 8;
         when "110011001001" => index <= 7;
         when "110011001010" => index <= 7;
         when "110011001011" => index <= 6;
         when "110011001100" => index <= 8;
         when "110011001101" => index <= 7;
         when "110011001110" => index <= 7;
         when "110011001111" => index <= 6;
         when "110011010000" => index <= 9;
         when "110011010001" => index <= 7;
         when "110011010010" => index <= 8;
         when "110011010011" => index <= 7;
         when "110011010100" => index <= 8;
         when "110011010101" => index <= 7;
         when "110011010110" => index <= 7;
         when "110011010111" => index <= 6;
         when "110011011000" => index <= 8;
         when "110011011001" => index <= 7;
         when "110011011010" => index <= 7;
         when "110011011011" => index <= 6;
         when "110011011100" => index <= 7;
         when "110011011101" => index <= 6;
         when "110011011110" => index <= 6;
         when "110011011111" => index <= 6;
         when "110011100000" => index <= 9;
         when "110011100001" => index <= 8;
         when "110011100010" => index <= 8;
         when "110011100011" => index <= 7;
         when "110011100100" => index <= 8;
         when "110011100101" => index <= 7;
         when "110011100110" => index <= 7;
         when "110011100111" => index <= 6;
         when "110011101000" => index <= 8;
         when "110011101001" => index <= 7;
         when "110011101010" => index <= 7;
         when "110011101011" => index <= 6;
         when "110011101100" => index <= 7;
         when "110011101101" => index <= 6;
         when "110011101110" => index <= 7;
         when "110011101111" => index <= 6;
         when "110011110000" => index <= 8;
         when "110011110001" => index <= 7;
         when "110011110010" => index <= 7;
         when "110011110011" => index <= 6;
         when "110011110100" => index <= 7;
         when "110011110101" => index <= 7;
         when "110011110110" => index <= 7;
         when "110011110111" => index <= 6;
         when "110011111000" => index <= 8;
         when "110011111001" => index <= 7;
         when "110011111010" => index <= 7;
         when "110011111011" => index <= 6;
         when "110011111100" => index <= 7;
         when "110011111101" => index <= 6;
         when "110011111110" => index <= 6;
         when "110011111111" => index <= 6;
         when "110100000000" => index <= 11;
         when "110100000001" => index <= 8;
         when "110100000010" => index <= 8;
         when "110100000011" => index <= 7;
         when "110100000100" => index <= 9;
         when "110100000101" => index <= 7;
         when "110100000110" => index <= 7;
         when "110100000111" => index <= 6;
         when "110100001000" => index <= 9;
         when "110100001001" => index <= 7;
         when "110100001010" => index <= 8;
         when "110100001011" => index <= 6;
         when "110100001100" => index <= 8;
         when "110100001101" => index <= 7;
         when "110100001110" => index <= 7;
         when "110100001111" => index <= 6;
         when "110100010000" => index <= 9;
         when "110100010001" => index <= 8;
         when "110100010010" => index <= 8;
         when "110100010011" => index <= 7;
         when "110100010100" => index <= 8;
         when "110100010101" => index <= 7;
         when "110100010110" => index <= 7;
         when "110100010111" => index <= 6;
         when "110100011000" => index <= 8;
         when "110100011001" => index <= 7;
         when "110100011010" => index <= 7;
         when "110100011011" => index <= 6;
         when "110100011100" => index <= 7;
         when "110100011101" => index <= 6;
         when "110100011110" => index <= 7;
         when "110100011111" => index <= 6;
         when "110100100000" => index <= 10;
         when "110100100001" => index <= 8;
         when "110100100010" => index <= 8;
         when "110100100011" => index <= 7;
         when "110100100100" => index <= 8;
         when "110100100101" => index <= 7;
         when "110100100110" => index <= 7;
         when "110100100111" => index <= 6;
         when "110100101000" => index <= 8;
         when "110100101001" => index <= 7;
         when "110100101010" => index <= 7;
         when "110100101011" => index <= 6;
         when "110100101100" => index <= 8;
         when "110100101101" => index <= 7;
         when "110100101110" => index <= 7;
         when "110100101111" => index <= 6;
         when "110100110000" => index <= 9;
         when "110100110001" => index <= 7;
         when "110100110010" => index <= 8;
         when "110100110011" => index <= 7;
         when "110100110100" => index <= 8;
         when "110100110101" => index <= 7;
         when "110100110110" => index <= 7;
         when "110100110111" => index <= 6;
         when "110100111000" => index <= 8;
         when "110100111001" => index <= 7;
         when "110100111010" => index <= 7;
         when "110100111011" => index <= 6;
         when "110100111100" => index <= 7;
         when "110100111101" => index <= 6;
         when "110100111110" => index <= 6;
         when "110100111111" => index <= 6;
         when "110101000000" => index <= 10;
         when "110101000001" => index <= 8;
         when "110101000010" => index <= 8;
         when "110101000011" => index <= 7;
         when "110101000100" => index <= 8;
         when "110101000101" => index <= 7;
         when "110101000110" => index <= 7;
         when "110101000111" => index <= 6;
         when "110101001000" => index <= 9;
         when "110101001001" => index <= 7;
         when "110101001010" => index <= 8;
         when "110101001011" => index <= 7;
         when "110101001100" => index <= 8;
         when "110101001101" => index <= 7;
         when "110101001110" => index <= 7;
         when "110101001111" => index <= 6;
         when "110101010000" => index <= 9;
         when "110101010001" => index <= 8;
         when "110101010010" => index <= 8;
         when "110101010011" => index <= 7;
         when "110101010100" => index <= 8;
         when "110101010101" => index <= 7;
         when "110101010110" => index <= 7;
         when "110101010111" => index <= 6;
         when "110101011000" => index <= 8;
         when "110101011001" => index <= 7;
         when "110101011010" => index <= 7;
         when "110101011011" => index <= 6;
         when "110101011100" => index <= 7;
         when "110101011101" => index <= 6;
         when "110101011110" => index <= 7;
         when "110101011111" => index <= 6;
         when "110101100000" => index <= 9;
         when "110101100001" => index <= 8;
         when "110101100010" => index <= 8;
         when "110101100011" => index <= 7;
         when "110101100100" => index <= 8;
         when "110101100101" => index <= 7;
         when "110101100110" => index <= 7;
         when "110101100111" => index <= 6;
         when "110101101000" => index <= 8;
         when "110101101001" => index <= 7;
         when "110101101010" => index <= 7;
         when "110101101011" => index <= 6;
         when "110101101100" => index <= 7;
         when "110101101101" => index <= 7;
         when "110101101110" => index <= 7;
         when "110101101111" => index <= 6;
         when "110101110000" => index <= 8;
         when "110101110001" => index <= 7;
         when "110101110010" => index <= 7;
         when "110101110011" => index <= 7;
         when "110101110100" => index <= 8;
         when "110101110101" => index <= 7;
         when "110101110110" => index <= 7;
         when "110101110111" => index <= 6;
         when "110101111000" => index <= 8;
         when "110101111001" => index <= 7;
         when "110101111010" => index <= 7;
         when "110101111011" => index <= 6;
         when "110101111100" => index <= 7;
         when "110101111101" => index <= 6;
         when "110101111110" => index <= 7;
         when "110101111111" => index <= 6;
         when "110110000000" => index <= 10;
         when "110110000001" => index <= 8;
         when "110110000010" => index <= 8;
         when "110110000011" => index <= 7;
         when "110110000100" => index <= 9;
         when "110110000101" => index <= 7;
         when "110110000110" => index <= 8;
         when "110110000111" => index <= 7;
         when "110110001000" => index <= 9;
         when "110110001001" => index <= 8;
         when "110110001010" => index <= 8;
         when "110110001011" => index <= 7;
         when "110110001100" => index <= 8;
         when "110110001101" => index <= 7;
         when "110110001110" => index <= 7;
         when "110110001111" => index <= 6;
         when "110110010000" => index <= 9;
         when "110110010001" => index <= 8;
         when "110110010010" => index <= 8;
         when "110110010011" => index <= 7;
         when "110110010100" => index <= 8;
         when "110110010101" => index <= 7;
         when "110110010110" => index <= 7;
         when "110110010111" => index <= 6;
         when "110110011000" => index <= 8;
         when "110110011001" => index <= 7;
         when "110110011010" => index <= 7;
         when "110110011011" => index <= 6;
         when "110110011100" => index <= 7;
         when "110110011101" => index <= 7;
         when "110110011110" => index <= 7;
         when "110110011111" => index <= 6;
         when "110110100000" => index <= 9;
         when "110110100001" => index <= 8;
         when "110110100010" => index <= 8;
         when "110110100011" => index <= 7;
         when "110110100100" => index <= 8;
         when "110110100101" => index <= 7;
         when "110110100110" => index <= 7;
         when "110110100111" => index <= 6;
         when "110110101000" => index <= 8;
         when "110110101001" => index <= 7;
         when "110110101010" => index <= 7;
         when "110110101011" => index <= 7;
         when "110110101100" => index <= 8;
         when "110110101101" => index <= 7;
         when "110110101110" => index <= 7;
         when "110110101111" => index <= 6;
         when "110110110000" => index <= 8;
         when "110110110001" => index <= 7;
         when "110110110010" => index <= 8;
         when "110110110011" => index <= 7;
         when "110110110100" => index <= 8;
         when "110110110101" => index <= 7;
         when "110110110110" => index <= 7;
         when "110110110111" => index <= 6;
         when "110110111000" => index <= 8;
         when "110110111001" => index <= 7;
         when "110110111010" => index <= 7;
         when "110110111011" => index <= 6;
         when "110110111100" => index <= 7;
         when "110110111101" => index <= 7;
         when "110110111110" => index <= 7;
         when "110110111111" => index <= 6;
         when "110111000000" => index <= 9;
         when "110111000001" => index <= 8;
         when "110111000010" => index <= 8;
         when "110111000011" => index <= 7;
         when "110111000100" => index <= 8;
         when "110111000101" => index <= 7;
         when "110111000110" => index <= 7;
         when "110111000111" => index <= 7;
         when "110111001000" => index <= 8;
         when "110111001001" => index <= 7;
         when "110111001010" => index <= 8;
         when "110111001011" => index <= 7;
         when "110111001100" => index <= 8;
         when "110111001101" => index <= 7;
         when "110111001110" => index <= 7;
         when "110111001111" => index <= 6;
         when "110111010000" => index <= 9;
         when "110111010001" => index <= 8;
         when "110111010010" => index <= 8;
         when "110111010011" => index <= 7;
         when "110111010100" => index <= 8;
         when "110111010101" => index <= 7;
         when "110111010110" => index <= 7;
         when "110111010111" => index <= 6;
         when "110111011000" => index <= 8;
         when "110111011001" => index <= 7;
         when "110111011010" => index <= 7;
         when "110111011011" => index <= 7;
         when "110111011100" => index <= 7;
         when "110111011101" => index <= 7;
         when "110111011110" => index <= 7;
         when "110111011111" => index <= 6;
         when "110111100000" => index <= 9;
         when "110111100001" => index <= 8;
         when "110111100010" => index <= 8;
         when "110111100011" => index <= 7;
         when "110111100100" => index <= 8;
         when "110111100101" => index <= 7;
         when "110111100110" => index <= 7;
         when "110111100111" => index <= 7;
         when "110111101000" => index <= 8;
         when "110111101001" => index <= 7;
         when "110111101010" => index <= 7;
         when "110111101011" => index <= 7;
         when "110111101100" => index <= 8;
         when "110111101101" => index <= 7;
         when "110111101110" => index <= 7;
         when "110111101111" => index <= 6;
         when "110111110000" => index <= 8;
         when "110111110001" => index <= 7;
         when "110111110010" => index <= 8;
         when "110111110011" => index <= 7;
         when "110111110100" => index <= 8;
         when "110111110101" => index <= 7;
         when "110111110110" => index <= 7;
         when "110111110111" => index <= 6;
         when "110111111000" => index <= 8;
         when "110111111001" => index <= 7;
         when "110111111010" => index <= 7;
         when "110111111011" => index <= 6;
         when "110111111100" => index <= 7;
         when "110111111101" => index <= 7;
         when "110111111110" => index <= 7;
         when "110111111111" => index <= 6;
         when "111000000000" => index <= 11;
         when "111000000001" => index <= 8;
         when "111000000010" => index <= 9;
         when "111000000011" => index <= 7;
         when "111000000100" => index <= 9;
         when "111000000101" => index <= 7;
         when "111000000110" => index <= 8;
         when "111000000111" => index <= 6;
         when "111000001000" => index <= 9;
         when "111000001001" => index <= 8;
         when "111000001010" => index <= 8;
         when "111000001011" => index <= 7;
         when "111000001100" => index <= 8;
         when "111000001101" => index <= 7;
         when "111000001110" => index <= 7;
         when "111000001111" => index <= 6;
         when "111000010000" => index <= 10;
         when "111000010001" => index <= 8;
         when "111000010010" => index <= 8;
         when "111000010011" => index <= 7;
         when "111000010100" => index <= 8;
         when "111000010101" => index <= 7;
         when "111000010110" => index <= 7;
         when "111000010111" => index <= 6;
         when "111000011000" => index <= 8;
         when "111000011001" => index <= 7;
         when "111000011010" => index <= 7;
         when "111000011011" => index <= 6;
         when "111000011100" => index <= 8;
         when "111000011101" => index <= 7;
         when "111000011110" => index <= 7;
         when "111000011111" => index <= 6;
         when "111000100000" => index <= 10;
         when "111000100001" => index <= 8;
         when "111000100010" => index <= 8;
         when "111000100011" => index <= 7;
         when "111000100100" => index <= 8;
         when "111000100101" => index <= 7;
         when "111000100110" => index <= 7;
         when "111000100111" => index <= 6;
         when "111000101000" => index <= 9;
         when "111000101001" => index <= 7;
         when "111000101010" => index <= 8;
         when "111000101011" => index <= 7;
         when "111000101100" => index <= 8;
         when "111000101101" => index <= 7;
         when "111000101110" => index <= 7;
         when "111000101111" => index <= 6;
         when "111000110000" => index <= 9;
         when "111000110001" => index <= 8;
         when "111000110010" => index <= 8;
         when "111000110011" => index <= 7;
         when "111000110100" => index <= 8;
         when "111000110101" => index <= 7;
         when "111000110110" => index <= 7;
         when "111000110111" => index <= 6;
         when "111000111000" => index <= 8;
         when "111000111001" => index <= 7;
         when "111000111010" => index <= 7;
         when "111000111011" => index <= 6;
         when "111000111100" => index <= 7;
         when "111000111101" => index <= 6;
         when "111000111110" => index <= 7;
         when "111000111111" => index <= 6;
         when "111001000000" => index <= 10;
         when "111001000001" => index <= 8;
         when "111001000010" => index <= 8;
         when "111001000011" => index <= 7;
         when "111001000100" => index <= 9;
         when "111001000101" => index <= 7;
         when "111001000110" => index <= 8;
         when "111001000111" => index <= 7;
         when "111001001000" => index <= 9;
         when "111001001001" => index <= 8;
         when "111001001010" => index <= 8;
         when "111001001011" => index <= 7;
         when "111001001100" => index <= 8;
         when "111001001101" => index <= 7;
         when "111001001110" => index <= 7;
         when "111001001111" => index <= 6;
         when "111001010000" => index <= 9;
         when "111001010001" => index <= 8;
         when "111001010010" => index <= 8;
         when "111001010011" => index <= 7;
         when "111001010100" => index <= 8;
         when "111001010101" => index <= 7;
         when "111001010110" => index <= 7;
         when "111001010111" => index <= 6;
         when "111001011000" => index <= 8;
         when "111001011001" => index <= 7;
         when "111001011010" => index <= 7;
         when "111001011011" => index <= 6;
         when "111001011100" => index <= 7;
         when "111001011101" => index <= 7;
         when "111001011110" => index <= 7;
         when "111001011111" => index <= 6;
         when "111001100000" => index <= 9;
         when "111001100001" => index <= 8;
         when "111001100010" => index <= 8;
         when "111001100011" => index <= 7;
         when "111001100100" => index <= 8;
         when "111001100101" => index <= 7;
         when "111001100110" => index <= 7;
         when "111001100111" => index <= 6;
         when "111001101000" => index <= 8;
         when "111001101001" => index <= 7;
         when "111001101010" => index <= 7;
         when "111001101011" => index <= 7;
         when "111001101100" => index <= 8;
         when "111001101101" => index <= 7;
         when "111001101110" => index <= 7;
         when "111001101111" => index <= 6;
         when "111001110000" => index <= 8;
         when "111001110001" => index <= 7;
         when "111001110010" => index <= 8;
         when "111001110011" => index <= 7;
         when "111001110100" => index <= 8;
         when "111001110101" => index <= 7;
         when "111001110110" => index <= 7;
         when "111001110111" => index <= 6;
         when "111001111000" => index <= 8;
         when "111001111001" => index <= 7;
         when "111001111010" => index <= 7;
         when "111001111011" => index <= 6;
         when "111001111100" => index <= 7;
         when "111001111101" => index <= 7;
         when "111001111110" => index <= 7;
         when "111001111111" => index <= 6;
         when "111010000000" => index <= 10;
         when "111010000001" => index <= 8;
         when "111010000010" => index <= 9;
         when "111010000011" => index <= 7;
         when "111010000100" => index <= 9;
         when "111010000101" => index <= 8;
         when "111010000110" => index <= 8;
         when "111010000111" => index <= 7;
         when "111010001000" => index <= 9;
         when "111010001001" => index <= 8;
         when "111010001010" => index <= 8;
         when "111010001011" => index <= 7;
         when "111010001100" => index <= 8;
         when "111010001101" => index <= 7;
         when "111010001110" => index <= 7;
         when "111010001111" => index <= 6;
         when "111010010000" => index <= 9;
         when "111010010001" => index <= 8;
         when "111010010010" => index <= 8;
         when "111010010011" => index <= 7;
         when "111010010100" => index <= 8;
         when "111010010101" => index <= 7;
         when "111010010110" => index <= 7;
         when "111010010111" => index <= 6;
         when "111010011000" => index <= 8;
         when "111010011001" => index <= 7;
         when "111010011010" => index <= 7;
         when "111010011011" => index <= 7;
         when "111010011100" => index <= 8;
         when "111010011101" => index <= 7;
         when "111010011110" => index <= 7;
         when "111010011111" => index <= 6;
         when "111010100000" => index <= 9;
         when "111010100001" => index <= 8;
         when "111010100010" => index <= 8;
         when "111010100011" => index <= 7;
         when "111010100100" => index <= 8;
         when "111010100101" => index <= 7;
         when "111010100110" => index <= 7;
         when "111010100111" => index <= 7;
         when "111010101000" => index <= 8;
         when "111010101001" => index <= 7;
         when "111010101010" => index <= 8;
         when "111010101011" => index <= 7;
         when "111010101100" => index <= 8;
         when "111010101101" => index <= 7;
         when "111010101110" => index <= 7;
         when "111010101111" => index <= 6;
         when "111010110000" => index <= 9;
         when "111010110001" => index <= 8;
         when "111010110010" => index <= 8;
         when "111010110011" => index <= 7;
         when "111010110100" => index <= 8;
         when "111010110101" => index <= 7;
         when "111010110110" => index <= 7;
         when "111010110111" => index <= 6;
         when "111010111000" => index <= 8;
         when "111010111001" => index <= 7;
         when "111010111010" => index <= 7;
         when "111010111011" => index <= 7;
         when "111010111100" => index <= 7;
         when "111010111101" => index <= 7;
         when "111010111110" => index <= 7;
         when "111010111111" => index <= 6;
         when "111011000000" => index <= 10;
         when "111011000001" => index <= 8;
         when "111011000010" => index <= 8;
         when "111011000011" => index <= 7;
         when "111011000100" => index <= 8;
         when "111011000101" => index <= 7;
         when "111011000110" => index <= 8;
         when "111011000111" => index <= 7;
         when "111011001000" => index <= 9;
         when "111011001001" => index <= 8;
         when "111011001010" => index <= 8;
         when "111011001011" => index <= 7;
         when "111011001100" => index <= 8;
         when "111011001101" => index <= 7;
         when "111011001110" => index <= 7;
         when "111011001111" => index <= 6;
         when "111011010000" => index <= 9;
         when "111011010001" => index <= 8;
         when "111011010010" => index <= 8;
         when "111011010011" => index <= 7;
         when "111011010100" => index <= 8;
         when "111011010101" => index <= 7;
         when "111011010110" => index <= 7;
         when "111011010111" => index <= 7;
         when "111011011000" => index <= 8;
         when "111011011001" => index <= 7;
         when "111011011010" => index <= 7;
         when "111011011011" => index <= 7;
         when "111011011100" => index <= 8;
         when "111011011101" => index <= 7;
         when "111011011110" => index <= 7;
         when "111011011111" => index <= 6;
         when "111011100000" => index <= 9;
         when "111011100001" => index <= 8;
         when "111011100010" => index <= 8;
         when "111011100011" => index <= 7;
         when "111011100100" => index <= 8;
         when "111011100101" => index <= 7;
         when "111011100110" => index <= 7;
         when "111011100111" => index <= 7;
         when "111011101000" => index <= 8;
         when "111011101001" => index <= 7;
         when "111011101010" => index <= 8;
         when "111011101011" => index <= 7;
         when "111011101100" => index <= 8;
         when "111011101101" => index <= 7;
         when "111011101110" => index <= 7;
         when "111011101111" => index <= 6;
         when "111011110000" => index <= 8;
         when "111011110001" => index <= 8;
         when "111011110010" => index <= 8;
         when "111011110011" => index <= 7;
         when "111011110100" => index <= 8;
         when "111011110101" => index <= 7;
         when "111011110110" => index <= 7;
         when "111011110111" => index <= 6;
         when "111011111000" => index <= 8;
         when "111011111001" => index <= 7;
         when "111011111010" => index <= 7;
         when "111011111011" => index <= 7;
         when "111011111100" => index <= 7;
         when "111011111101" => index <= 7;
         when "111011111110" => index <= 7;
         when "111011111111" => index <= 6;
         when "111100000000" => index <= 10;
         when "111100000001" => index <= 9;
         when "111100000010" => index <= 9;
         when "111100000011" => index <= 8;
         when "111100000100" => index <= 9;
         when "111100000101" => index <= 8;
         when "111100000110" => index <= 8;
         when "111100000111" => index <= 7;
         when "111100001000" => index <= 9;
         when "111100001001" => index <= 8;
         when "111100001010" => index <= 8;
         when "111100001011" => index <= 7;
         when "111100001100" => index <= 8;
         when "111100001101" => index <= 7;
         when "111100001110" => index <= 7;
         when "111100001111" => index <= 6;
         when "111100010000" => index <= 9;
         when "111100010001" => index <= 8;
         when "111100010010" => index <= 8;
         when "111100010011" => index <= 7;
         when "111100010100" => index <= 8;
         when "111100010101" => index <= 7;
         when "111100010110" => index <= 7;
         when "111100010111" => index <= 7;
         when "111100011000" => index <= 8;
         when "111100011001" => index <= 7;
         when "111100011010" => index <= 8;
         when "111100011011" => index <= 7;
         when "111100011100" => index <= 8;
         when "111100011101" => index <= 7;
         when "111100011110" => index <= 7;
         when "111100011111" => index <= 6;
         when "111100100000" => index <= 10;
         when "111100100001" => index <= 8;
         when "111100100010" => index <= 8;
         when "111100100011" => index <= 7;
         when "111100100100" => index <= 8;
         when "111100100101" => index <= 7;
         when "111100100110" => index <= 8;
         when "111100100111" => index <= 7;
         when "111100101000" => index <= 9;
         when "111100101001" => index <= 8;
         when "111100101010" => index <= 8;
         when "111100101011" => index <= 7;
         when "111100101100" => index <= 8;
         when "111100101101" => index <= 7;
         when "111100101110" => index <= 7;
         when "111100101111" => index <= 6;
         when "111100110000" => index <= 9;
         when "111100110001" => index <= 8;
         when "111100110010" => index <= 8;
         when "111100110011" => index <= 7;
         when "111100110100" => index <= 8;
         when "111100110101" => index <= 7;
         when "111100110110" => index <= 7;
         when "111100110111" => index <= 7;
         when "111100111000" => index <= 8;
         when "111100111001" => index <= 7;
         when "111100111010" => index <= 7;
         when "111100111011" => index <= 7;
         when "111100111100" => index <= 8;
         when "111100111101" => index <= 7;
         when "111100111110" => index <= 7;
         when "111100111111" => index <= 6;
         when "111101000000" => index <= 10;
         when "111101000001" => index <= 8;
         when "111101000010" => index <= 8;
         when "111101000011" => index <= 7;
         when "111101000100" => index <= 9;
         when "111101000101" => index <= 8;
         when "111101000110" => index <= 8;
         when "111101000111" => index <= 7;
         when "111101001000" => index <= 9;
         when "111101001001" => index <= 8;
         when "111101001010" => index <= 8;
         when "111101001011" => index <= 7;
         when "111101001100" => index <= 8;
         when "111101001101" => index <= 7;
         when "111101001110" => index <= 7;
         when "111101001111" => index <= 7;
         when "111101010000" => index <= 9;
         when "111101010001" => index <= 8;
         when "111101010010" => index <= 8;
         when "111101010011" => index <= 7;
         when "111101010100" => index <= 8;
         when "111101010101" => index <= 7;
         when "111101010110" => index <= 7;
         when "111101010111" => index <= 7;
         when "111101011000" => index <= 8;
         when "111101011001" => index <= 7;
         when "111101011010" => index <= 8;
         when "111101011011" => index <= 7;
         when "111101011100" => index <= 8;
         when "111101011101" => index <= 7;
         when "111101011110" => index <= 7;
         when "111101011111" => index <= 6;
         when "111101100000" => index <= 9;
         when "111101100001" => index <= 8;
         when "111101100010" => index <= 8;
         when "111101100011" => index <= 7;
         when "111101100100" => index <= 8;
         when "111101100101" => index <= 7;
         when "111101100110" => index <= 8;
         when "111101100111" => index <= 7;
         when "111101101000" => index <= 8;
         when "111101101001" => index <= 8;
         when "111101101010" => index <= 8;
         when "111101101011" => index <= 7;
         when "111101101100" => index <= 8;
         when "111101101101" => index <= 7;
         when "111101101110" => index <= 7;
         when "111101101111" => index <= 6;
         when "111101110000" => index <= 9;
         when "111101110001" => index <= 8;
         when "111101110010" => index <= 8;
         when "111101110011" => index <= 7;
         when "111101110100" => index <= 8;
         when "111101110101" => index <= 7;
         when "111101110110" => index <= 7;
         when "111101110111" => index <= 7;
         when "111101111000" => index <= 8;
         when "111101111001" => index <= 7;
         when "111101111010" => index <= 7;
         when "111101111011" => index <= 7;
         when "111101111100" => index <= 7;
         when "111101111101" => index <= 7;
         when "111101111110" => index <= 7;
         when "111101111111" => index <= 6;
         when "111110000000" => index <= 10;
         when "111110000001" => index <= 8;
         when "111110000010" => index <= 9;
         when "111110000011" => index <= 8;
         when "111110000100" => index <= 9;
         when "111110000101" => index <= 8;
         when "111110000110" => index <= 8;
         when "111110000111" => index <= 7;
         when "111110001000" => index <= 9;
         when "111110001001" => index <= 8;
         when "111110001010" => index <= 8;
         when "111110001011" => index <= 7;
         when "111110001100" => index <= 8;
         when "111110001101" => index <= 7;
         when "111110001110" => index <= 7;
         when "111110001111" => index <= 7;
         when "111110010000" => index <= 9;
         when "111110010001" => index <= 8;
         when "111110010010" => index <= 8;
         when "111110010011" => index <= 7;
         when "111110010100" => index <= 8;
         when "111110010101" => index <= 7;
         when "111110010110" => index <= 8;
         when "111110010111" => index <= 7;
         when "111110011000" => index <= 8;
         when "111110011001" => index <= 8;
         when "111110011010" => index <= 8;
         when "111110011011" => index <= 7;
         when "111110011100" => index <= 8;
         when "111110011101" => index <= 7;
         when "111110011110" => index <= 7;
         when "111110011111" => index <= 6;
         when "111110100000" => index <= 9;
         when "111110100001" => index <= 8;
         when "111110100010" => index <= 8;
         when "111110100011" => index <= 7;
         when "111110100100" => index <= 8;
         when "111110100101" => index <= 8;
         when "111110100110" => index <= 8;
         when "111110100111" => index <= 7;
         when "111110101000" => index <= 9;
         when "111110101001" => index <= 8;
         when "111110101010" => index <= 8;
         when "111110101011" => index <= 7;
         when "111110101100" => index <= 8;
         when "111110101101" => index <= 7;
         when "111110101110" => index <= 7;
         when "111110101111" => index <= 7;
         when "111110110000" => index <= 9;
         when "111110110001" => index <= 8;
         when "111110110010" => index <= 8;
         when "111110110011" => index <= 7;
         when "111110110100" => index <= 8;
         when "111110110101" => index <= 7;
         when "111110110110" => index <= 7;
         when "111110110111" => index <= 7;
         when "111110111000" => index <= 8;
         when "111110111001" => index <= 7;
         when "111110111010" => index <= 7;
         when "111110111011" => index <= 7;
         when "111110111100" => index <= 8;
         when "111110111101" => index <= 7;
         when "111110111110" => index <= 7;
         when "111110111111" => index <= 6;
         when "111111000000" => index <= 10;
         when "111111000001" => index <= 8;
         when "111111000010" => index <= 8;
         when "111111000011" => index <= 8;
         when "111111000100" => index <= 9;
         when "111111000101" => index <= 8;
         when "111111000110" => index <= 8;
         when "111111000111" => index <= 7;
         when "111111001000" => index <= 9;
         when "111111001001" => index <= 8;
         when "111111001010" => index <= 8;
         when "111111001011" => index <= 7;
         when "111111001100" => index <= 8;
         when "111111001101" => index <= 7;
         when "111111001110" => index <= 7;
         when "111111001111" => index <= 7;
         when "111111010000" => index <= 9;
         when "111111010001" => index <= 8;
         when "111111010010" => index <= 8;
         when "111111010011" => index <= 7;
         when "111111010100" => index <= 8;
         when "111111010101" => index <= 7;
         when "111111010110" => index <= 7;
         when "111111010111" => index <= 7;
         when "111111011000" => index <= 8;
         when "111111011001" => index <= 7;
         when "111111011010" => index <= 8;
         when "111111011011" => index <= 7;
         when "111111011100" => index <= 8;
         when "111111011101" => index <= 7;
         when "111111011110" => index <= 7;
         when "111111011111" => index <= 7;
         when "111111100000" => index <= 9;
         when "111111100001" => index <= 8;
         when "111111100010" => index <= 8;
         when "111111100011" => index <= 7;
         when "111111100100" => index <= 8;
         when "111111100101" => index <= 7;
         when "111111100110" => index <= 8;
         when "111111100111" => index <= 7;
         when "111111101000" => index <= 8;
         when "111111101001" => index <= 8;
         when "111111101010" => index <= 8;
         when "111111101011" => index <= 7;
         when "111111101100" => index <= 8;
         when "111111101101" => index <= 7;
         when "111111101110" => index <= 7;
         when "111111101111" => index <= 7;
         when "111111110000" => index <= 8;
         when "111111110001" => index <= 8;
         when "111111110010" => index <= 8;
         when "111111110011" => index <= 7;
         when "111111110100" => index <= 8;
         when "111111110101" => index <= 7;
         when "111111110110" => index <= 7;
         when "111111110111" => index <= 7;
         when "111111111000" => index <= 8;
         when "111111111001" => index <= 7;
         when "111111111010" => index <= 7;
         when "111111111011" => index <= 7;
         when "111111111100" => index <= 8;
         when "111111111101" => index <= 7;
         when "111111111110" => index <= 7;
         when "111111111111" => index <= 6;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;


  gen_13 : if (length = 13) generate
  begin
    process (clk) is
    begin
      if (rising_edge(clk)) then
        case din is
         when "0000000000000" => index <= 0;
         when "0000000000001" => index <= 1;
         when "0000000000010" => index <= 2;
         when "0000000000011" => index <= 2;
         when "0000000000100" => index <= 3;
         when "0000000000101" => index <= 2;
         when "0000000000110" => index <= 2;
         when "0000000000111" => index <= 2;
         when "0000000001000" => index <= 4;
         when "0000000001001" => index <= 2;
         when "0000000001010" => index <= 3;
         when "0000000001011" => index <= 2;
         when "0000000001100" => index <= 4;
         when "0000000001101" => index <= 3;
         when "0000000001110" => index <= 3;
         when "0000000001111" => index <= 2;
         when "0000000010000" => index <= 5;
         when "0000000010001" => index <= 3;
         when "0000000010010" => index <= 4;
         when "0000000010011" => index <= 3;
         when "0000000010100" => index <= 4;
         when "0000000010101" => index <= 3;
         when "0000000010110" => index <= 3;
         when "0000000010111" => index <= 3;
         when "0000000011000" => index <= 4;
         when "0000000011001" => index <= 3;
         when "0000000011010" => index <= 4;
         when "0000000011011" => index <= 3;
         when "0000000011100" => index <= 4;
         when "0000000011101" => index <= 3;
         when "0000000011110" => index <= 4;
         when "0000000011111" => index <= 3;
         when "0000000100000" => index <= 6;
         when "0000000100001" => index <= 4;
         when "0000000100010" => index <= 4;
         when "0000000100011" => index <= 3;
         when "0000000100100" => index <= 4;
         when "0000000100101" => index <= 3;
         when "0000000100110" => index <= 4;
         when "0000000100111" => index <= 3;
         when "0000000101000" => index <= 5;
         when "0000000101001" => index <= 4;
         when "0000000101010" => index <= 4;
         when "0000000101011" => index <= 3;
         when "0000000101100" => index <= 4;
         when "0000000101101" => index <= 4;
         when "0000000101110" => index <= 4;
         when "0000000101111" => index <= 3;
         when "0000000110000" => index <= 6;
         when "0000000110001" => index <= 4;
         when "0000000110010" => index <= 4;
         when "0000000110011" => index <= 4;
         when "0000000110100" => index <= 5;
         when "0000000110101" => index <= 4;
         when "0000000110110" => index <= 4;
         when "0000000110111" => index <= 3;
         when "0000000111000" => index <= 5;
         when "0000000111001" => index <= 4;
         when "0000000111010" => index <= 4;
         when "0000000111011" => index <= 4;
         when "0000000111100" => index <= 4;
         when "0000000111101" => index <= 4;
         when "0000000111110" => index <= 4;
         when "0000000111111" => index <= 4;
         when "0000001000000" => index <= 7;
         when "0000001000001" => index <= 4;
         when "0000001000010" => index <= 4;
         when "0000001000011" => index <= 3;
         when "0000001000100" => index <= 5;
         when "0000001000101" => index <= 4;
         when "0000001000110" => index <= 4;
         when "0000001000111" => index <= 3;
         when "0000001001000" => index <= 6;
         when "0000001001001" => index <= 4;
         when "0000001001010" => index <= 4;
         when "0000001001011" => index <= 4;
         when "0000001001100" => index <= 5;
         when "0000001001101" => index <= 4;
         when "0000001001110" => index <= 4;
         when "0000001001111" => index <= 3;
         when "0000001010000" => index <= 6;
         when "0000001010001" => index <= 4;
         when "0000001010010" => index <= 5;
         when "0000001010011" => index <= 4;
         when "0000001010100" => index <= 5;
         when "0000001010101" => index <= 4;
         when "0000001010110" => index <= 4;
         when "0000001010111" => index <= 4;
         when "0000001011000" => index <= 5;
         when "0000001011001" => index <= 4;
         when "0000001011010" => index <= 4;
         when "0000001011011" => index <= 4;
         when "0000001011100" => index <= 5;
         when "0000001011101" => index <= 4;
         when "0000001011110" => index <= 4;
         when "0000001011111" => index <= 4;
         when "0000001100000" => index <= 6;
         when "0000001100001" => index <= 5;
         when "0000001100010" => index <= 5;
         when "0000001100011" => index <= 4;
         when "0000001100100" => index <= 5;
         when "0000001100101" => index <= 4;
         when "0000001100110" => index <= 4;
         when "0000001100111" => index <= 4;
         when "0000001101000" => index <= 6;
         when "0000001101001" => index <= 4;
         when "0000001101010" => index <= 5;
         when "0000001101011" => index <= 4;
         when "0000001101100" => index <= 5;
         when "0000001101101" => index <= 4;
         when "0000001101110" => index <= 4;
         when "0000001101111" => index <= 4;
         when "0000001110000" => index <= 6;
         when "0000001110001" => index <= 5;
         when "0000001110010" => index <= 5;
         when "0000001110011" => index <= 4;
         when "0000001110100" => index <= 5;
         when "0000001110101" => index <= 4;
         when "0000001110110" => index <= 5;
         when "0000001110111" => index <= 4;
         when "0000001111000" => index <= 6;
         when "0000001111001" => index <= 5;
         when "0000001111010" => index <= 5;
         when "0000001111011" => index <= 4;
         when "0000001111100" => index <= 5;
         when "0000001111101" => index <= 4;
         when "0000001111110" => index <= 4;
         when "0000001111111" => index <= 4;
         when "0000010000000" => index <= 8;
         when "0000010000001" => index <= 4;
         when "0000010000010" => index <= 5;
         when "0000010000011" => index <= 4;
         when "0000010000100" => index <= 6;
         when "0000010000101" => index <= 4;
         when "0000010000110" => index <= 4;
         when "0000010000111" => index <= 4;
         when "0000010001000" => index <= 6;
         when "0000010001001" => index <= 4;
         when "0000010001010" => index <= 5;
         when "0000010001011" => index <= 4;
         when "0000010001100" => index <= 5;
         when "0000010001101" => index <= 4;
         when "0000010001110" => index <= 4;
         when "0000010001111" => index <= 4;
         when "0000010010000" => index <= 6;
         when "0000010010001" => index <= 5;
         when "0000010010010" => index <= 5;
         when "0000010010011" => index <= 4;
         when "0000010010100" => index <= 5;
         when "0000010010101" => index <= 4;
         when "0000010010110" => index <= 4;
         when "0000010010111" => index <= 4;
         when "0000010011000" => index <= 6;
         when "0000010011001" => index <= 4;
         when "0000010011010" => index <= 5;
         when "0000010011011" => index <= 4;
         when "0000010011100" => index <= 5;
         when "0000010011101" => index <= 4;
         when "0000010011110" => index <= 4;
         when "0000010011111" => index <= 4;
         when "0000010100000" => index <= 7;
         when "0000010100001" => index <= 5;
         when "0000010100010" => index <= 5;
         when "0000010100011" => index <= 4;
         when "0000010100100" => index <= 6;
         when "0000010100101" => index <= 4;
         when "0000010100110" => index <= 5;
         when "0000010100111" => index <= 4;
         when "0000010101000" => index <= 6;
         when "0000010101001" => index <= 5;
         when "0000010101010" => index <= 5;
         when "0000010101011" => index <= 4;
         when "0000010101100" => index <= 5;
         when "0000010101101" => index <= 4;
         when "0000010101110" => index <= 5;
         when "0000010101111" => index <= 4;
         when "0000010110000" => index <= 6;
         when "0000010110001" => index <= 5;
         when "0000010110010" => index <= 5;
         when "0000010110011" => index <= 4;
         when "0000010110100" => index <= 6;
         when "0000010110101" => index <= 5;
         when "0000010110110" => index <= 5;
         when "0000010110111" => index <= 4;
         when "0000010111000" => index <= 6;
         when "0000010111001" => index <= 5;
         when "0000010111010" => index <= 5;
         when "0000010111011" => index <= 4;
         when "0000010111100" => index <= 5;
         when "0000010111101" => index <= 4;
         when "0000010111110" => index <= 5;
         when "0000010111111" => index <= 4;
         when "0000011000000" => index <= 8;
         when "0000011000001" => index <= 5;
         when "0000011000010" => index <= 6;
         when "0000011000011" => index <= 4;
         when "0000011000100" => index <= 6;
         when "0000011000101" => index <= 5;
         when "0000011000110" => index <= 5;
         when "0000011000111" => index <= 4;
         when "0000011001000" => index <= 6;
         when "0000011001001" => index <= 5;
         when "0000011001010" => index <= 5;
         when "0000011001011" => index <= 4;
         when "0000011001100" => index <= 6;
         when "0000011001101" => index <= 5;
         when "0000011001110" => index <= 5;
         when "0000011001111" => index <= 4;
         when "0000011010000" => index <= 7;
         when "0000011010001" => index <= 5;
         when "0000011010010" => index <= 6;
         when "0000011010011" => index <= 5;
         when "0000011010100" => index <= 6;
         when "0000011010101" => index <= 5;
         when "0000011010110" => index <= 5;
         when "0000011010111" => index <= 4;
         when "0000011011000" => index <= 6;
         when "0000011011001" => index <= 5;
         when "0000011011010" => index <= 5;
         when "0000011011011" => index <= 4;
         when "0000011011100" => index <= 5;
         when "0000011011101" => index <= 5;
         when "0000011011110" => index <= 5;
         when "0000011011111" => index <= 4;
         when "0000011100000" => index <= 7;
         when "0000011100001" => index <= 6;
         when "0000011100010" => index <= 6;
         when "0000011100011" => index <= 5;
         when "0000011100100" => index <= 6;
         when "0000011100101" => index <= 5;
         when "0000011100110" => index <= 5;
         when "0000011100111" => index <= 4;
         when "0000011101000" => index <= 6;
         when "0000011101001" => index <= 5;
         when "0000011101010" => index <= 5;
         when "0000011101011" => index <= 5;
         when "0000011101100" => index <= 6;
         when "0000011101101" => index <= 5;
         when "0000011101110" => index <= 5;
         when "0000011101111" => index <= 4;
         when "0000011110000" => index <= 6;
         when "0000011110001" => index <= 5;
         when "0000011110010" => index <= 6;
         when "0000011110011" => index <= 5;
         when "0000011110100" => index <= 6;
         when "0000011110101" => index <= 5;
         when "0000011110110" => index <= 5;
         when "0000011110111" => index <= 5;
         when "0000011111000" => index <= 6;
         when "0000011111001" => index <= 5;
         when "0000011111010" => index <= 5;
         when "0000011111011" => index <= 5;
         when "0000011111100" => index <= 6;
         when "0000011111101" => index <= 5;
         when "0000011111110" => index <= 5;
         when "0000011111111" => index <= 4;
         when "0000100000000" => index <= 9;
         when "0000100000001" => index <= 5;
         when "0000100000010" => index <= 6;
         when "0000100000011" => index <= 4;
         when "0000100000100" => index <= 6;
         when "0000100000101" => index <= 4;
         when "0000100000110" => index <= 5;
         when "0000100000111" => index <= 4;
         when "0000100001000" => index <= 6;
         when "0000100001001" => index <= 5;
         when "0000100001010" => index <= 5;
         when "0000100001011" => index <= 4;
         when "0000100001100" => index <= 5;
         when "0000100001101" => index <= 4;
         when "0000100001110" => index <= 4;
         when "0000100001111" => index <= 4;
         when "0000100010000" => index <= 7;
         when "0000100010001" => index <= 5;
         when "0000100010010" => index <= 5;
         when "0000100010011" => index <= 4;
         when "0000100010100" => index <= 6;
         when "0000100010101" => index <= 4;
         when "0000100010110" => index <= 5;
         when "0000100010111" => index <= 4;
         when "0000100011000" => index <= 6;
         when "0000100011001" => index <= 5;
         when "0000100011010" => index <= 5;
         when "0000100011011" => index <= 4;
         when "0000100011100" => index <= 5;
         when "0000100011101" => index <= 4;
         when "0000100011110" => index <= 5;
         when "0000100011111" => index <= 4;
         when "0000100100000" => index <= 8;
         when "0000100100001" => index <= 5;
         when "0000100100010" => index <= 6;
         when "0000100100011" => index <= 4;
         when "0000100100100" => index <= 6;
         when "0000100100101" => index <= 5;
         when "0000100100110" => index <= 5;
         when "0000100100111" => index <= 4;
         when "0000100101000" => index <= 6;
         when "0000100101001" => index <= 5;
         when "0000100101010" => index <= 5;
         when "0000100101011" => index <= 4;
         when "0000100101100" => index <= 6;
         when "0000100101101" => index <= 5;
         when "0000100101110" => index <= 5;
         when "0000100101111" => index <= 4;
         when "0000100110000" => index <= 7;
         when "0000100110001" => index <= 5;
         when "0000100110010" => index <= 6;
         when "0000100110011" => index <= 5;
         when "0000100110100" => index <= 6;
         when "0000100110101" => index <= 5;
         when "0000100110110" => index <= 5;
         when "0000100110111" => index <= 4;
         when "0000100111000" => index <= 6;
         when "0000100111001" => index <= 5;
         when "0000100111010" => index <= 5;
         when "0000100111011" => index <= 4;
         when "0000100111100" => index <= 5;
         when "0000100111101" => index <= 5;
         when "0000100111110" => index <= 5;
         when "0000100111111" => index <= 4;
         when "0000101000000" => index <= 8;
         when "0000101000001" => index <= 6;
         when "0000101000010" => index <= 6;
         when "0000101000011" => index <= 5;
         when "0000101000100" => index <= 6;
         when "0000101000101" => index <= 5;
         when "0000101000110" => index <= 5;
         when "0000101000111" => index <= 4;
         when "0000101001000" => index <= 7;
         when "0000101001001" => index <= 5;
         when "0000101001010" => index <= 6;
         when "0000101001011" => index <= 5;
         when "0000101001100" => index <= 6;
         when "0000101001101" => index <= 5;
         when "0000101001110" => index <= 5;
         when "0000101001111" => index <= 4;
         when "0000101010000" => index <= 7;
         when "0000101010001" => index <= 6;
         when "0000101010010" => index <= 6;
         when "0000101010011" => index <= 5;
         when "0000101010100" => index <= 6;
         when "0000101010101" => index <= 5;
         when "0000101010110" => index <= 5;
         when "0000101010111" => index <= 4;
         when "0000101011000" => index <= 6;
         when "0000101011001" => index <= 5;
         when "0000101011010" => index <= 5;
         when "0000101011011" => index <= 5;
         when "0000101011100" => index <= 6;
         when "0000101011101" => index <= 5;
         when "0000101011110" => index <= 5;
         when "0000101011111" => index <= 4;
         when "0000101100000" => index <= 7;
         when "0000101100001" => index <= 6;
         when "0000101100010" => index <= 6;
         when "0000101100011" => index <= 5;
         when "0000101100100" => index <= 6;
         when "0000101100101" => index <= 5;
         when "0000101100110" => index <= 5;
         when "0000101100111" => index <= 5;
         when "0000101101000" => index <= 6;
         when "0000101101001" => index <= 5;
         when "0000101101010" => index <= 6;
         when "0000101101011" => index <= 5;
         when "0000101101100" => index <= 6;
         when "0000101101101" => index <= 5;
         when "0000101101110" => index <= 5;
         when "0000101101111" => index <= 5;
         when "0000101110000" => index <= 7;
         when "0000101110001" => index <= 6;
         when "0000101110010" => index <= 6;
         when "0000101110011" => index <= 5;
         when "0000101110100" => index <= 6;
         when "0000101110101" => index <= 5;
         when "0000101110110" => index <= 5;
         when "0000101110111" => index <= 5;
         when "0000101111000" => index <= 6;
         when "0000101111001" => index <= 5;
         when "0000101111010" => index <= 6;
         when "0000101111011" => index <= 5;
         when "0000101111100" => index <= 6;
         when "0000101111101" => index <= 5;
         when "0000101111110" => index <= 5;
         when "0000101111111" => index <= 5;
         when "0000110000000" => index <= 8;
         when "0000110000001" => index <= 6;
         when "0000110000010" => index <= 6;
         when "0000110000011" => index <= 5;
         when "0000110000100" => index <= 7;
         when "0000110000101" => index <= 5;
         when "0000110000110" => index <= 6;
         when "0000110000111" => index <= 5;
         when "0000110001000" => index <= 7;
         when "0000110001001" => index <= 6;
         when "0000110001010" => index <= 6;
         when "0000110001011" => index <= 5;
         when "0000110001100" => index <= 6;
         when "0000110001101" => index <= 5;
         when "0000110001110" => index <= 5;
         when "0000110001111" => index <= 4;
         when "0000110010000" => index <= 7;
         when "0000110010001" => index <= 6;
         when "0000110010010" => index <= 6;
         when "0000110010011" => index <= 5;
         when "0000110010100" => index <= 6;
         when "0000110010101" => index <= 5;
         when "0000110010110" => index <= 5;
         when "0000110010111" => index <= 5;
         when "0000110011000" => index <= 6;
         when "0000110011001" => index <= 5;
         when "0000110011010" => index <= 6;
         when "0000110011011" => index <= 5;
         when "0000110011100" => index <= 6;
         when "0000110011101" => index <= 5;
         when "0000110011110" => index <= 5;
         when "0000110011111" => index <= 5;
         when "0000110100000" => index <= 8;
         when "0000110100001" => index <= 6;
         when "0000110100010" => index <= 6;
         when "0000110100011" => index <= 5;
         when "0000110100100" => index <= 6;
         when "0000110100101" => index <= 5;
         when "0000110100110" => index <= 6;
         when "0000110100111" => index <= 5;
         when "0000110101000" => index <= 7;
         when "0000110101001" => index <= 6;
         when "0000110101010" => index <= 6;
         when "0000110101011" => index <= 5;
         when "0000110101100" => index <= 6;
         when "0000110101101" => index <= 5;
         when "0000110101110" => index <= 5;
         when "0000110101111" => index <= 5;
         when "0000110110000" => index <= 7;
         when "0000110110001" => index <= 6;
         when "0000110110010" => index <= 6;
         when "0000110110011" => index <= 5;
         when "0000110110100" => index <= 6;
         when "0000110110101" => index <= 5;
         when "0000110110110" => index <= 6;
         when "0000110110111" => index <= 5;
         when "0000110111000" => index <= 6;
         when "0000110111001" => index <= 6;
         when "0000110111010" => index <= 6;
         when "0000110111011" => index <= 5;
         when "0000110111100" => index <= 6;
         when "0000110111101" => index <= 5;
         when "0000110111110" => index <= 5;
         when "0000110111111" => index <= 5;
         when "0000111000000" => index <= 8;
         when "0000111000001" => index <= 6;
         when "0000111000010" => index <= 6;
         when "0000111000011" => index <= 5;
         when "0000111000100" => index <= 7;
         when "0000111000101" => index <= 6;
         when "0000111000110" => index <= 6;
         when "0000111000111" => index <= 5;
         when "0000111001000" => index <= 7;
         when "0000111001001" => index <= 6;
         when "0000111001010" => index <= 6;
         when "0000111001011" => index <= 5;
         when "0000111001100" => index <= 6;
         when "0000111001101" => index <= 5;
         when "0000111001110" => index <= 6;
         when "0000111001111" => index <= 5;
         when "0000111010000" => index <= 7;
         when "0000111010001" => index <= 6;
         when "0000111010010" => index <= 6;
         when "0000111010011" => index <= 5;
         when "0000111010100" => index <= 6;
         when "0000111010101" => index <= 6;
         when "0000111010110" => index <= 6;
         when "0000111010111" => index <= 5;
         when "0000111011000" => index <= 7;
         when "0000111011001" => index <= 6;
         when "0000111011010" => index <= 6;
         when "0000111011011" => index <= 5;
         when "0000111011100" => index <= 6;
         when "0000111011101" => index <= 5;
         when "0000111011110" => index <= 5;
         when "0000111011111" => index <= 5;
         when "0000111100000" => index <= 8;
         when "0000111100001" => index <= 6;
         when "0000111100010" => index <= 6;
         when "0000111100011" => index <= 6;
         when "0000111100100" => index <= 7;
         when "0000111100101" => index <= 6;
         when "0000111100110" => index <= 6;
         when "0000111100111" => index <= 5;
         when "0000111101000" => index <= 7;
         when "0000111101001" => index <= 6;
         when "0000111101010" => index <= 6;
         when "0000111101011" => index <= 5;
         when "0000111101100" => index <= 6;
         when "0000111101101" => index <= 5;
         when "0000111101110" => index <= 6;
         when "0000111101111" => index <= 5;
         when "0000111110000" => index <= 7;
         when "0000111110001" => index <= 6;
         when "0000111110010" => index <= 6;
         when "0000111110011" => index <= 5;
         when "0000111110100" => index <= 6;
         when "0000111110101" => index <= 6;
         when "0000111110110" => index <= 6;
         when "0000111110111" => index <= 5;
         when "0000111111000" => index <= 6;
         when "0000111111001" => index <= 6;
         when "0000111111010" => index <= 6;
         when "0000111111011" => index <= 5;
         when "0000111111100" => index <= 6;
         when "0000111111101" => index <= 5;
         when "0000111111110" => index <= 6;
         when "0000111111111" => index <= 5;
         when "0001000000000" => index <= 10;
         when "0001000000001" => index <= 6;
         when "0001000000010" => index <= 6;
         when "0001000000011" => index <= 4;
         when "0001000000100" => index <= 6;
         when "0001000000101" => index <= 5;
         when "0001000000110" => index <= 5;
         when "0001000000111" => index <= 4;
         when "0001000001000" => index <= 7;
         when "0001000001001" => index <= 5;
         when "0001000001010" => index <= 5;
         when "0001000001011" => index <= 4;
         when "0001000001100" => index <= 6;
         when "0001000001101" => index <= 4;
         when "0001000001110" => index <= 5;
         when "0001000001111" => index <= 4;
         when "0001000010000" => index <= 8;
         when "0001000010001" => index <= 5;
         when "0001000010010" => index <= 6;
         when "0001000010011" => index <= 4;
         when "0001000010100" => index <= 6;
         when "0001000010101" => index <= 5;
         when "0001000010110" => index <= 5;
         when "0001000010111" => index <= 4;
         when "0001000011000" => index <= 6;
         when "0001000011001" => index <= 5;
         when "0001000011010" => index <= 5;
         when "0001000011011" => index <= 4;
         when "0001000011100" => index <= 6;
         when "0001000011101" => index <= 5;
         when "0001000011110" => index <= 5;
         when "0001000011111" => index <= 4;
         when "0001000100000" => index <= 8;
         when "0001000100001" => index <= 6;
         when "0001000100010" => index <= 6;
         when "0001000100011" => index <= 5;
         when "0001000100100" => index <= 6;
         when "0001000100101" => index <= 5;
         when "0001000100110" => index <= 5;
         when "0001000100111" => index <= 4;
         when "0001000101000" => index <= 7;
         when "0001000101001" => index <= 5;
         when "0001000101010" => index <= 6;
         when "0001000101011" => index <= 5;
         when "0001000101100" => index <= 6;
         when "0001000101101" => index <= 5;
         when "0001000101110" => index <= 5;
         when "0001000101111" => index <= 4;
         when "0001000110000" => index <= 7;
         when "0001000110001" => index <= 6;
         when "0001000110010" => index <= 6;
         when "0001000110011" => index <= 5;
         when "0001000110100" => index <= 6;
         when "0001000110101" => index <= 5;
         when "0001000110110" => index <= 5;
         when "0001000110111" => index <= 4;
         when "0001000111000" => index <= 6;
         when "0001000111001" => index <= 5;
         when "0001000111010" => index <= 5;
         when "0001000111011" => index <= 5;
         when "0001000111100" => index <= 6;
         when "0001000111101" => index <= 5;
         when "0001000111110" => index <= 5;
         when "0001000111111" => index <= 4;
         when "0001001000000" => index <= 8;
         when "0001001000001" => index <= 6;
         when "0001001000010" => index <= 6;
         when "0001001000011" => index <= 5;
         when "0001001000100" => index <= 7;
         when "0001001000101" => index <= 5;
         when "0001001000110" => index <= 6;
         when "0001001000111" => index <= 5;
         when "0001001001000" => index <= 7;
         when "0001001001001" => index <= 6;
         when "0001001001010" => index <= 6;
         when "0001001001011" => index <= 5;
         when "0001001001100" => index <= 6;
         when "0001001001101" => index <= 5;
         when "0001001001110" => index <= 5;
         when "0001001001111" => index <= 4;
         when "0001001010000" => index <= 7;
         when "0001001010001" => index <= 6;
         when "0001001010010" => index <= 6;
         when "0001001010011" => index <= 5;
         when "0001001010100" => index <= 6;
         when "0001001010101" => index <= 5;
         when "0001001010110" => index <= 5;
         when "0001001010111" => index <= 5;
         when "0001001011000" => index <= 6;
         when "0001001011001" => index <= 5;
         when "0001001011010" => index <= 6;
         when "0001001011011" => index <= 5;
         when "0001001011100" => index <= 6;
         when "0001001011101" => index <= 5;
         when "0001001011110" => index <= 5;
         when "0001001011111" => index <= 5;
         when "0001001100000" => index <= 8;
         when "0001001100001" => index <= 6;
         when "0001001100010" => index <= 6;
         when "0001001100011" => index <= 5;
         when "0001001100100" => index <= 6;
         when "0001001100101" => index <= 5;
         when "0001001100110" => index <= 6;
         when "0001001100111" => index <= 5;
         when "0001001101000" => index <= 7;
         when "0001001101001" => index <= 6;
         when "0001001101010" => index <= 6;
         when "0001001101011" => index <= 5;
         when "0001001101100" => index <= 6;
         when "0001001101101" => index <= 5;
         when "0001001101110" => index <= 5;
         when "0001001101111" => index <= 5;
         when "0001001110000" => index <= 7;
         when "0001001110001" => index <= 6;
         when "0001001110010" => index <= 6;
         when "0001001110011" => index <= 5;
         when "0001001110100" => index <= 6;
         when "0001001110101" => index <= 5;
         when "0001001110110" => index <= 6;
         when "0001001110111" => index <= 5;
         when "0001001111000" => index <= 6;
         when "0001001111001" => index <= 6;
         when "0001001111010" => index <= 6;
         when "0001001111011" => index <= 5;
         when "0001001111100" => index <= 6;
         when "0001001111101" => index <= 5;
         when "0001001111110" => index <= 5;
         when "0001001111111" => index <= 5;
         when "0001010000000" => index <= 9;
         when "0001010000001" => index <= 6;
         when "0001010000010" => index <= 7;
         when "0001010000011" => index <= 5;
         when "0001010000100" => index <= 7;
         when "0001010000101" => index <= 6;
         when "0001010000110" => index <= 6;
         when "0001010000111" => index <= 5;
         when "0001010001000" => index <= 7;
         when "0001010001001" => index <= 6;
         when "0001010001010" => index <= 6;
         when "0001010001011" => index <= 5;
         when "0001010001100" => index <= 6;
         when "0001010001101" => index <= 5;
         when "0001010001110" => index <= 5;
         when "0001010001111" => index <= 5;
         when "0001010010000" => index <= 8;
         when "0001010010001" => index <= 6;
         when "0001010010010" => index <= 6;
         when "0001010010011" => index <= 5;
         when "0001010010100" => index <= 6;
         when "0001010010101" => index <= 5;
         when "0001010010110" => index <= 6;
         when "0001010010111" => index <= 5;
         when "0001010011000" => index <= 7;
         when "0001010011001" => index <= 6;
         when "0001010011010" => index <= 6;
         when "0001010011011" => index <= 5;
         when "0001010011100" => index <= 6;
         when "0001010011101" => index <= 5;
         when "0001010011110" => index <= 5;
         when "0001010011111" => index <= 5;
         when "0001010100000" => index <= 8;
         when "0001010100001" => index <= 6;
         when "0001010100010" => index <= 6;
         when "0001010100011" => index <= 5;
         when "0001010100100" => index <= 7;
         when "0001010100101" => index <= 6;
         when "0001010100110" => index <= 6;
         when "0001010100111" => index <= 5;
         when "0001010101000" => index <= 7;
         when "0001010101001" => index <= 6;
         when "0001010101010" => index <= 6;
         when "0001010101011" => index <= 5;
         when "0001010101100" => index <= 6;
         when "0001010101101" => index <= 5;
         when "0001010101110" => index <= 6;
         when "0001010101111" => index <= 5;
         when "0001010110000" => index <= 7;
         when "0001010110001" => index <= 6;
         when "0001010110010" => index <= 6;
         when "0001010110011" => index <= 5;
         when "0001010110100" => index <= 6;
         when "0001010110101" => index <= 6;
         when "0001010110110" => index <= 6;
         when "0001010110111" => index <= 5;
         when "0001010111000" => index <= 7;
         when "0001010111001" => index <= 6;
         when "0001010111010" => index <= 6;
         when "0001010111011" => index <= 5;
         when "0001010111100" => index <= 6;
         when "0001010111101" => index <= 5;
         when "0001010111110" => index <= 5;
         when "0001010111111" => index <= 5;
         when "0001011000000" => index <= 8;
         when "0001011000001" => index <= 6;
         when "0001011000010" => index <= 7;
         when "0001011000011" => index <= 6;
         when "0001011000100" => index <= 7;
         when "0001011000101" => index <= 6;
         when "0001011000110" => index <= 6;
         when "0001011000111" => index <= 5;
         when "0001011001000" => index <= 7;
         when "0001011001001" => index <= 6;
         when "0001011001010" => index <= 6;
         when "0001011001011" => index <= 5;
         when "0001011001100" => index <= 6;
         when "0001011001101" => index <= 6;
         when "0001011001110" => index <= 6;
         when "0001011001111" => index <= 5;
         when "0001011010000" => index <= 8;
         when "0001011010001" => index <= 6;
         when "0001011010010" => index <= 6;
         when "0001011010011" => index <= 6;
         when "0001011010100" => index <= 7;
         when "0001011010101" => index <= 6;
         when "0001011010110" => index <= 6;
         when "0001011010111" => index <= 5;
         when "0001011011000" => index <= 7;
         when "0001011011001" => index <= 6;
         when "0001011011010" => index <= 6;
         when "0001011011011" => index <= 5;
         when "0001011011100" => index <= 6;
         when "0001011011101" => index <= 5;
         when "0001011011110" => index <= 6;
         when "0001011011111" => index <= 5;
         when "0001011100000" => index <= 8;
         when "0001011100001" => index <= 6;
         when "0001011100010" => index <= 7;
         when "0001011100011" => index <= 6;
         when "0001011100100" => index <= 7;
         when "0001011100101" => index <= 6;
         when "0001011100110" => index <= 6;
         when "0001011100111" => index <= 5;
         when "0001011101000" => index <= 7;
         when "0001011101001" => index <= 6;
         when "0001011101010" => index <= 6;
         when "0001011101011" => index <= 5;
         when "0001011101100" => index <= 6;
         when "0001011101101" => index <= 6;
         when "0001011101110" => index <= 6;
         when "0001011101111" => index <= 5;
         when "0001011110000" => index <= 7;
         when "0001011110001" => index <= 6;
         when "0001011110010" => index <= 6;
         when "0001011110011" => index <= 6;
         when "0001011110100" => index <= 6;
         when "0001011110101" => index <= 6;
         when "0001011110110" => index <= 6;
         when "0001011110111" => index <= 5;
         when "0001011111000" => index <= 7;
         when "0001011111001" => index <= 6;
         when "0001011111010" => index <= 6;
         when "0001011111011" => index <= 5;
         when "0001011111100" => index <= 6;
         when "0001011111101" => index <= 6;
         when "0001011111110" => index <= 6;
         when "0001011111111" => index <= 5;
         when "0001100000000" => index <= 10;
         when "0001100000001" => index <= 7;
         when "0001100000010" => index <= 7;
         when "0001100000011" => index <= 6;
         when "0001100000100" => index <= 7;
         when "0001100000101" => index <= 6;
         when "0001100000110" => index <= 6;
         when "0001100000111" => index <= 5;
         when "0001100001000" => index <= 8;
         when "0001100001001" => index <= 6;
         when "0001100001010" => index <= 6;
         when "0001100001011" => index <= 5;
         when "0001100001100" => index <= 6;
         when "0001100001101" => index <= 5;
         when "0001100001110" => index <= 6;
         when "0001100001111" => index <= 5;
         when "0001100010000" => index <= 8;
         when "0001100010001" => index <= 6;
         when "0001100010010" => index <= 6;
         when "0001100010011" => index <= 5;
         when "0001100010100" => index <= 7;
         when "0001100010101" => index <= 6;
         when "0001100010110" => index <= 6;
         when "0001100010111" => index <= 5;
         when "0001100011000" => index <= 7;
         when "0001100011001" => index <= 6;
         when "0001100011010" => index <= 6;
         when "0001100011011" => index <= 5;
         when "0001100011100" => index <= 6;
         when "0001100011101" => index <= 5;
         when "0001100011110" => index <= 6;
         when "0001100011111" => index <= 5;
         when "0001100100000" => index <= 8;
         when "0001100100001" => index <= 6;
         when "0001100100010" => index <= 7;
         when "0001100100011" => index <= 6;
         when "0001100100100" => index <= 7;
         when "0001100100101" => index <= 6;
         when "0001100100110" => index <= 6;
         when "0001100100111" => index <= 5;
         when "0001100101000" => index <= 7;
         when "0001100101001" => index <= 6;
         when "0001100101010" => index <= 6;
         when "0001100101011" => index <= 5;
         when "0001100101100" => index <= 6;
         when "0001100101101" => index <= 6;
         when "0001100101110" => index <= 6;
         when "0001100101111" => index <= 5;
         when "0001100110000" => index <= 8;
         when "0001100110001" => index <= 6;
         when "0001100110010" => index <= 6;
         when "0001100110011" => index <= 6;
         when "0001100110100" => index <= 7;
         when "0001100110101" => index <= 6;
         when "0001100110110" => index <= 6;
         when "0001100110111" => index <= 5;
         when "0001100111000" => index <= 7;
         when "0001100111001" => index <= 6;
         when "0001100111010" => index <= 6;
         when "0001100111011" => index <= 5;
         when "0001100111100" => index <= 6;
         when "0001100111101" => index <= 5;
         when "0001100111110" => index <= 6;
         when "0001100111111" => index <= 5;
         when "0001101000000" => index <= 9;
         when "0001101000001" => index <= 7;
         when "0001101000010" => index <= 7;
         when "0001101000011" => index <= 6;
         when "0001101000100" => index <= 7;
         when "0001101000101" => index <= 6;
         when "0001101000110" => index <= 6;
         when "0001101000111" => index <= 5;
         when "0001101001000" => index <= 8;
         when "0001101001001" => index <= 6;
         when "0001101001010" => index <= 6;
         when "0001101001011" => index <= 6;
         when "0001101001100" => index <= 7;
         when "0001101001101" => index <= 6;
         when "0001101001110" => index <= 6;
         when "0001101001111" => index <= 5;
         when "0001101010000" => index <= 8;
         when "0001101010001" => index <= 6;
         when "0001101010010" => index <= 7;
         when "0001101010011" => index <= 6;
         when "0001101010100" => index <= 7;
         when "0001101010101" => index <= 6;
         when "0001101010110" => index <= 6;
         when "0001101010111" => index <= 5;
         when "0001101011000" => index <= 7;
         when "0001101011001" => index <= 6;
         when "0001101011010" => index <= 6;
         when "0001101011011" => index <= 5;
         when "0001101011100" => index <= 6;
         when "0001101011101" => index <= 6;
         when "0001101011110" => index <= 6;
         when "0001101011111" => index <= 5;
         when "0001101100000" => index <= 8;
         when "0001101100001" => index <= 7;
         when "0001101100010" => index <= 7;
         when "0001101100011" => index <= 6;
         when "0001101100100" => index <= 7;
         when "0001101100101" => index <= 6;
         when "0001101100110" => index <= 6;
         when "0001101100111" => index <= 5;
         when "0001101101000" => index <= 7;
         when "0001101101001" => index <= 6;
         when "0001101101010" => index <= 6;
         when "0001101101011" => index <= 6;
         when "0001101101100" => index <= 6;
         when "0001101101101" => index <= 6;
         when "0001101101110" => index <= 6;
         when "0001101101111" => index <= 5;
         when "0001101110000" => index <= 7;
         when "0001101110001" => index <= 6;
         when "0001101110010" => index <= 6;
         when "0001101110011" => index <= 6;
         when "0001101110100" => index <= 7;
         when "0001101110101" => index <= 6;
         when "0001101110110" => index <= 6;
         when "0001101110111" => index <= 5;
         when "0001101111000" => index <= 7;
         when "0001101111001" => index <= 6;
         when "0001101111010" => index <= 6;
         when "0001101111011" => index <= 6;
         when "0001101111100" => index <= 6;
         when "0001101111101" => index <= 6;
         when "0001101111110" => index <= 6;
         when "0001101111111" => index <= 5;
         when "0001110000000" => index <= 9;
         when "0001110000001" => index <= 7;
         when "0001110000010" => index <= 7;
         when "0001110000011" => index <= 6;
         when "0001110000100" => index <= 8;
         when "0001110000101" => index <= 6;
         when "0001110000110" => index <= 6;
         when "0001110000111" => index <= 6;
         when "0001110001000" => index <= 8;
         when "0001110001001" => index <= 6;
         when "0001110001010" => index <= 7;
         when "0001110001011" => index <= 6;
         when "0001110001100" => index <= 7;
         when "0001110001101" => index <= 6;
         when "0001110001110" => index <= 6;
         when "0001110001111" => index <= 5;
         when "0001110010000" => index <= 8;
         when "0001110010001" => index <= 7;
         when "0001110010010" => index <= 7;
         when "0001110010011" => index <= 6;
         when "0001110010100" => index <= 7;
         when "0001110010101" => index <= 6;
         when "0001110010110" => index <= 6;
         when "0001110010111" => index <= 5;
         when "0001110011000" => index <= 7;
         when "0001110011001" => index <= 6;
         when "0001110011010" => index <= 6;
         when "0001110011011" => index <= 6;
         when "0001110011100" => index <= 6;
         when "0001110011101" => index <= 6;
         when "0001110011110" => index <= 6;
         when "0001110011111" => index <= 5;
         when "0001110100000" => index <= 8;
         when "0001110100001" => index <= 7;
         when "0001110100010" => index <= 7;
         when "0001110100011" => index <= 6;
         when "0001110100100" => index <= 7;
         when "0001110100101" => index <= 6;
         when "0001110100110" => index <= 6;
         when "0001110100111" => index <= 6;
         when "0001110101000" => index <= 7;
         when "0001110101001" => index <= 6;
         when "0001110101010" => index <= 6;
         when "0001110101011" => index <= 6;
         when "0001110101100" => index <= 7;
         when "0001110101101" => index <= 6;
         when "0001110101110" => index <= 6;
         when "0001110101111" => index <= 5;
         when "0001110110000" => index <= 8;
         when "0001110110001" => index <= 6;
         when "0001110110010" => index <= 7;
         when "0001110110011" => index <= 6;
         when "0001110110100" => index <= 7;
         when "0001110110101" => index <= 6;
         when "0001110110110" => index <= 6;
         when "0001110110111" => index <= 6;
         when "0001110111000" => index <= 7;
         when "0001110111001" => index <= 6;
         when "0001110111010" => index <= 6;
         when "0001110111011" => index <= 6;
         when "0001110111100" => index <= 6;
         when "0001110111101" => index <= 6;
         when "0001110111110" => index <= 6;
         when "0001110111111" => index <= 5;
         when "0001111000000" => index <= 8;
         when "0001111000001" => index <= 7;
         when "0001111000010" => index <= 7;
         when "0001111000011" => index <= 6;
         when "0001111000100" => index <= 7;
         when "0001111000101" => index <= 6;
         when "0001111000110" => index <= 6;
         when "0001111000111" => index <= 6;
         when "0001111001000" => index <= 8;
         when "0001111001001" => index <= 6;
         when "0001111001010" => index <= 7;
         when "0001111001011" => index <= 6;
         when "0001111001100" => index <= 7;
         when "0001111001101" => index <= 6;
         when "0001111001110" => index <= 6;
         when "0001111001111" => index <= 6;
         when "0001111010000" => index <= 8;
         when "0001111010001" => index <= 7;
         when "0001111010010" => index <= 7;
         when "0001111010011" => index <= 6;
         when "0001111010100" => index <= 7;
         when "0001111010101" => index <= 6;
         when "0001111010110" => index <= 6;
         when "0001111010111" => index <= 6;
         when "0001111011000" => index <= 7;
         when "0001111011001" => index <= 6;
         when "0001111011010" => index <= 6;
         when "0001111011011" => index <= 6;
         when "0001111011100" => index <= 7;
         when "0001111011101" => index <= 6;
         when "0001111011110" => index <= 6;
         when "0001111011111" => index <= 5;
         when "0001111100000" => index <= 8;
         when "0001111100001" => index <= 7;
         when "0001111100010" => index <= 7;
         when "0001111100011" => index <= 6;
         when "0001111100100" => index <= 7;
         when "0001111100101" => index <= 6;
         when "0001111100110" => index <= 6;
         when "0001111100111" => index <= 6;
         when "0001111101000" => index <= 7;
         when "0001111101001" => index <= 6;
         when "0001111101010" => index <= 7;
         when "0001111101011" => index <= 6;
         when "0001111101100" => index <= 7;
         when "0001111101101" => index <= 6;
         when "0001111101110" => index <= 6;
         when "0001111101111" => index <= 6;
         when "0001111110000" => index <= 8;
         when "0001111110001" => index <= 7;
         when "0001111110010" => index <= 7;
         when "0001111110011" => index <= 6;
         when "0001111110100" => index <= 7;
         when "0001111110101" => index <= 6;
         when "0001111110110" => index <= 6;
         when "0001111110111" => index <= 6;
         when "0001111111000" => index <= 7;
         when "0001111111001" => index <= 6;
         when "0001111111010" => index <= 6;
         when "0001111111011" => index <= 6;
         when "0001111111100" => index <= 6;
         when "0001111111101" => index <= 6;
         when "0001111111110" => index <= 6;
         when "0001111111111" => index <= 6;
         when "0010000000000" => index <= 11;
         when "0010000000001" => index <= 6;
         when "0010000000010" => index <= 6;
         when "0010000000011" => index <= 5;
         when "0010000000100" => index <= 7;
         when "0010000000101" => index <= 5;
         when "0010000000110" => index <= 5;
         when "0010000000111" => index <= 4;
         when "0010000001000" => index <= 8;
         when "0010000001001" => index <= 5;
         when "0010000001010" => index <= 6;
         when "0010000001011" => index <= 4;
         when "0010000001100" => index <= 6;
         when "0010000001101" => index <= 5;
         when "0010000001110" => index <= 5;
         when "0010000001111" => index <= 4;
         when "0010000010000" => index <= 8;
         when "0010000010001" => index <= 6;
         when "0010000010010" => index <= 6;
         when "0010000010011" => index <= 5;
         when "0010000010100" => index <= 6;
         when "0010000010101" => index <= 5;
         when "0010000010110" => index <= 5;
         when "0010000010111" => index <= 4;
         when "0010000011000" => index <= 7;
         when "0010000011001" => index <= 5;
         when "0010000011010" => index <= 6;
         when "0010000011011" => index <= 5;
         when "0010000011100" => index <= 6;
         when "0010000011101" => index <= 5;
         when "0010000011110" => index <= 5;
         when "0010000011111" => index <= 4;
         when "0010000100000" => index <= 8;
         when "0010000100001" => index <= 6;
         when "0010000100010" => index <= 6;
         when "0010000100011" => index <= 5;
         when "0010000100100" => index <= 7;
         when "0010000100101" => index <= 5;
         when "0010000100110" => index <= 6;
         when "0010000100111" => index <= 5;
         when "0010000101000" => index <= 7;
         when "0010000101001" => index <= 6;
         when "0010000101010" => index <= 6;
         when "0010000101011" => index <= 5;
         when "0010000101100" => index <= 6;
         when "0010000101101" => index <= 5;
         when "0010000101110" => index <= 5;
         when "0010000101111" => index <= 4;
         when "0010000110000" => index <= 7;
         when "0010000110001" => index <= 6;
         when "0010000110010" => index <= 6;
         when "0010000110011" => index <= 5;
         when "0010000110100" => index <= 6;
         when "0010000110101" => index <= 5;
         when "0010000110110" => index <= 5;
         when "0010000110111" => index <= 5;
         when "0010000111000" => index <= 6;
         when "0010000111001" => index <= 5;
         when "0010000111010" => index <= 6;
         when "0010000111011" => index <= 5;
         when "0010000111100" => index <= 6;
         when "0010000111101" => index <= 5;
         when "0010000111110" => index <= 5;
         when "0010000111111" => index <= 5;
         when "0010001000000" => index <= 9;
         when "0010001000001" => index <= 6;
         when "0010001000010" => index <= 7;
         when "0010001000011" => index <= 5;
         when "0010001000100" => index <= 7;
         when "0010001000101" => index <= 6;
         when "0010001000110" => index <= 6;
         when "0010001000111" => index <= 5;
         when "0010001001000" => index <= 7;
         when "0010001001001" => index <= 6;
         when "0010001001010" => index <= 6;
         when "0010001001011" => index <= 5;
         when "0010001001100" => index <= 6;
         when "0010001001101" => index <= 5;
         when "0010001001110" => index <= 5;
         when "0010001001111" => index <= 5;
         when "0010001010000" => index <= 8;
         when "0010001010001" => index <= 6;
         when "0010001010010" => index <= 6;
         when "0010001010011" => index <= 5;
         when "0010001010100" => index <= 6;
         when "0010001010101" => index <= 5;
         when "0010001010110" => index <= 6;
         when "0010001010111" => index <= 5;
         when "0010001011000" => index <= 7;
         when "0010001011001" => index <= 6;
         when "0010001011010" => index <= 6;
         when "0010001011011" => index <= 5;
         when "0010001011100" => index <= 6;
         when "0010001011101" => index <= 5;
         when "0010001011110" => index <= 5;
         when "0010001011111" => index <= 5;
         when "0010001100000" => index <= 8;
         when "0010001100001" => index <= 6;
         when "0010001100010" => index <= 6;
         when "0010001100011" => index <= 5;
         when "0010001100100" => index <= 7;
         when "0010001100101" => index <= 6;
         when "0010001100110" => index <= 6;
         when "0010001100111" => index <= 5;
         when "0010001101000" => index <= 7;
         when "0010001101001" => index <= 6;
         when "0010001101010" => index <= 6;
         when "0010001101011" => index <= 5;
         when "0010001101100" => index <= 6;
         when "0010001101101" => index <= 5;
         when "0010001101110" => index <= 6;
         when "0010001101111" => index <= 5;
         when "0010001110000" => index <= 7;
         when "0010001110001" => index <= 6;
         when "0010001110010" => index <= 6;
         when "0010001110011" => index <= 5;
         when "0010001110100" => index <= 6;
         when "0010001110101" => index <= 6;
         when "0010001110110" => index <= 6;
         when "0010001110111" => index <= 5;
         when "0010001111000" => index <= 7;
         when "0010001111001" => index <= 6;
         when "0010001111010" => index <= 6;
         when "0010001111011" => index <= 5;
         when "0010001111100" => index <= 6;
         when "0010001111101" => index <= 5;
         when "0010001111110" => index <= 5;
         when "0010001111111" => index <= 5;
         when "0010010000000" => index <= 10;
         when "0010010000001" => index <= 7;
         when "0010010000010" => index <= 7;
         when "0010010000011" => index <= 6;
         when "0010010000100" => index <= 7;
         when "0010010000101" => index <= 6;
         when "0010010000110" => index <= 6;
         when "0010010000111" => index <= 5;
         when "0010010001000" => index <= 8;
         when "0010010001001" => index <= 6;
         when "0010010001010" => index <= 6;
         when "0010010001011" => index <= 5;
         when "0010010001100" => index <= 6;
         when "0010010001101" => index <= 5;
         when "0010010001110" => index <= 6;
         when "0010010001111" => index <= 5;
         when "0010010010000" => index <= 8;
         when "0010010010001" => index <= 6;
         when "0010010010010" => index <= 6;
         when "0010010010011" => index <= 5;
         when "0010010010100" => index <= 7;
         when "0010010010101" => index <= 6;
         when "0010010010110" => index <= 6;
         when "0010010010111" => index <= 5;
         when "0010010011000" => index <= 7;
         when "0010010011001" => index <= 6;
         when "0010010011010" => index <= 6;
         when "0010010011011" => index <= 5;
         when "0010010011100" => index <= 6;
         when "0010010011101" => index <= 5;
         when "0010010011110" => index <= 6;
         when "0010010011111" => index <= 5;
         when "0010010100000" => index <= 8;
         when "0010010100001" => index <= 6;
         when "0010010100010" => index <= 7;
         when "0010010100011" => index <= 6;
         when "0010010100100" => index <= 7;
         when "0010010100101" => index <= 6;
         when "0010010100110" => index <= 6;
         when "0010010100111" => index <= 5;
         when "0010010101000" => index <= 7;
         when "0010010101001" => index <= 6;
         when "0010010101010" => index <= 6;
         when "0010010101011" => index <= 5;
         when "0010010101100" => index <= 6;
         when "0010010101101" => index <= 6;
         when "0010010101110" => index <= 6;
         when "0010010101111" => index <= 5;
         when "0010010110000" => index <= 8;
         when "0010010110001" => index <= 6;
         when "0010010110010" => index <= 6;
         when "0010010110011" => index <= 6;
         when "0010010110100" => index <= 7;
         when "0010010110101" => index <= 6;
         when "0010010110110" => index <= 6;
         when "0010010110111" => index <= 5;
         when "0010010111000" => index <= 7;
         when "0010010111001" => index <= 6;
         when "0010010111010" => index <= 6;
         when "0010010111011" => index <= 5;
         when "0010010111100" => index <= 6;
         when "0010010111101" => index <= 5;
         when "0010010111110" => index <= 6;
         when "0010010111111" => index <= 5;
         when "0010011000000" => index <= 9;
         when "0010011000001" => index <= 7;
         when "0010011000010" => index <= 7;
         when "0010011000011" => index <= 6;
         when "0010011000100" => index <= 7;
         when "0010011000101" => index <= 6;
         when "0010011000110" => index <= 6;
         when "0010011000111" => index <= 5;
         when "0010011001000" => index <= 8;
         when "0010011001001" => index <= 6;
         when "0010011001010" => index <= 6;
         when "0010011001011" => index <= 6;
         when "0010011001100" => index <= 7;
         when "0010011001101" => index <= 6;
         when "0010011001110" => index <= 6;
         when "0010011001111" => index <= 5;
         when "0010011010000" => index <= 8;
         when "0010011010001" => index <= 6;
         when "0010011010010" => index <= 7;
         when "0010011010011" => index <= 6;
         when "0010011010100" => index <= 7;
         when "0010011010101" => index <= 6;
         when "0010011010110" => index <= 6;
         when "0010011010111" => index <= 5;
         when "0010011011000" => index <= 7;
         when "0010011011001" => index <= 6;
         when "0010011011010" => index <= 6;
         when "0010011011011" => index <= 5;
         when "0010011011100" => index <= 6;
         when "0010011011101" => index <= 6;
         when "0010011011110" => index <= 6;
         when "0010011011111" => index <= 5;
         when "0010011100000" => index <= 8;
         when "0010011100001" => index <= 7;
         when "0010011100010" => index <= 7;
         when "0010011100011" => index <= 6;
         when "0010011100100" => index <= 7;
         when "0010011100101" => index <= 6;
         when "0010011100110" => index <= 6;
         when "0010011100111" => index <= 5;
         when "0010011101000" => index <= 7;
         when "0010011101001" => index <= 6;
         when "0010011101010" => index <= 6;
         when "0010011101011" => index <= 6;
         when "0010011101100" => index <= 6;
         when "0010011101101" => index <= 6;
         when "0010011101110" => index <= 6;
         when "0010011101111" => index <= 5;
         when "0010011110000" => index <= 7;
         when "0010011110001" => index <= 6;
         when "0010011110010" => index <= 6;
         when "0010011110011" => index <= 6;
         when "0010011110100" => index <= 7;
         when "0010011110101" => index <= 6;
         when "0010011110110" => index <= 6;
         when "0010011110111" => index <= 5;
         when "0010011111000" => index <= 7;
         when "0010011111001" => index <= 6;
         when "0010011111010" => index <= 6;
         when "0010011111011" => index <= 6;
         when "0010011111100" => index <= 6;
         when "0010011111101" => index <= 6;
         when "0010011111110" => index <= 6;
         when "0010011111111" => index <= 5;
         when "0010100000000" => index <= 10;
         when "0010100000001" => index <= 7;
         when "0010100000010" => index <= 7;
         when "0010100000011" => index <= 6;
         when "0010100000100" => index <= 8;
         when "0010100000101" => index <= 6;
         when "0010100000110" => index <= 6;
         when "0010100000111" => index <= 5;
         when "0010100001000" => index <= 8;
         when "0010100001001" => index <= 6;
         when "0010100001010" => index <= 6;
         when "0010100001011" => index <= 5;
         when "0010100001100" => index <= 7;
         when "0010100001101" => index <= 6;
         when "0010100001110" => index <= 6;
         when "0010100001111" => index <= 5;
         when "0010100010000" => index <= 8;
         when "0010100010001" => index <= 6;
         when "0010100010010" => index <= 7;
         when "0010100010011" => index <= 6;
         when "0010100010100" => index <= 7;
         when "0010100010101" => index <= 6;
         when "0010100010110" => index <= 6;
         when "0010100010111" => index <= 5;
         when "0010100011000" => index <= 7;
         when "0010100011001" => index <= 6;
         when "0010100011010" => index <= 6;
         when "0010100011011" => index <= 5;
         when "0010100011100" => index <= 6;
         when "0010100011101" => index <= 6;
         when "0010100011110" => index <= 6;
         when "0010100011111" => index <= 5;
         when "0010100100000" => index <= 9;
         when "0010100100001" => index <= 7;
         when "0010100100010" => index <= 7;
         when "0010100100011" => index <= 6;
         when "0010100100100" => index <= 7;
         when "0010100100101" => index <= 6;
         when "0010100100110" => index <= 6;
         when "0010100100111" => index <= 5;
         when "0010100101000" => index <= 8;
         when "0010100101001" => index <= 6;
         when "0010100101010" => index <= 6;
         when "0010100101011" => index <= 6;
         when "0010100101100" => index <= 7;
         when "0010100101101" => index <= 6;
         when "0010100101110" => index <= 6;
         when "0010100101111" => index <= 5;
         when "0010100110000" => index <= 8;
         when "0010100110001" => index <= 6;
         when "0010100110010" => index <= 7;
         when "0010100110011" => index <= 6;
         when "0010100110100" => index <= 7;
         when "0010100110101" => index <= 6;
         when "0010100110110" => index <= 6;
         when "0010100110111" => index <= 5;
         when "0010100111000" => index <= 7;
         when "0010100111001" => index <= 6;
         when "0010100111010" => index <= 6;
         when "0010100111011" => index <= 5;
         when "0010100111100" => index <= 6;
         when "0010100111101" => index <= 6;
         when "0010100111110" => index <= 6;
         when "0010100111111" => index <= 5;
         when "0010101000000" => index <= 9;
         when "0010101000001" => index <= 7;
         when "0010101000010" => index <= 7;
         when "0010101000011" => index <= 6;
         when "0010101000100" => index <= 8;
         when "0010101000101" => index <= 6;
         when "0010101000110" => index <= 6;
         when "0010101000111" => index <= 6;
         when "0010101001000" => index <= 8;
         when "0010101001001" => index <= 6;
         when "0010101001010" => index <= 7;
         when "0010101001011" => index <= 6;
         when "0010101001100" => index <= 7;
         when "0010101001101" => index <= 6;
         when "0010101001110" => index <= 6;
         when "0010101001111" => index <= 5;
         when "0010101010000" => index <= 8;
         when "0010101010001" => index <= 7;
         when "0010101010010" => index <= 7;
         when "0010101010011" => index <= 6;
         when "0010101010100" => index <= 7;
         when "0010101010101" => index <= 6;
         when "0010101010110" => index <= 6;
         when "0010101010111" => index <= 5;
         when "0010101011000" => index <= 7;
         when "0010101011001" => index <= 6;
         when "0010101011010" => index <= 6;
         when "0010101011011" => index <= 6;
         when "0010101011100" => index <= 6;
         when "0010101011101" => index <= 6;
         when "0010101011110" => index <= 6;
         when "0010101011111" => index <= 5;
         when "0010101100000" => index <= 8;
         when "0010101100001" => index <= 7;
         when "0010101100010" => index <= 7;
         when "0010101100011" => index <= 6;
         when "0010101100100" => index <= 7;
         when "0010101100101" => index <= 6;
         when "0010101100110" => index <= 6;
         when "0010101100111" => index <= 6;
         when "0010101101000" => index <= 7;
         when "0010101101001" => index <= 6;
         when "0010101101010" => index <= 6;
         when "0010101101011" => index <= 6;
         when "0010101101100" => index <= 7;
         when "0010101101101" => index <= 6;
         when "0010101101110" => index <= 6;
         when "0010101101111" => index <= 5;
         when "0010101110000" => index <= 8;
         when "0010101110001" => index <= 6;
         when "0010101110010" => index <= 7;
         when "0010101110011" => index <= 6;
         when "0010101110100" => index <= 7;
         when "0010101110101" => index <= 6;
         when "0010101110110" => index <= 6;
         when "0010101110111" => index <= 6;
         when "0010101111000" => index <= 7;
         when "0010101111001" => index <= 6;
         when "0010101111010" => index <= 6;
         when "0010101111011" => index <= 6;
         when "0010101111100" => index <= 6;
         when "0010101111101" => index <= 6;
         when "0010101111110" => index <= 6;
         when "0010101111111" => index <= 5;
         when "0010110000000" => index <= 9;
         when "0010110000001" => index <= 7;
         when "0010110000010" => index <= 8;
         when "0010110000011" => index <= 6;
         when "0010110000100" => index <= 8;
         when "0010110000101" => index <= 6;
         when "0010110000110" => index <= 7;
         when "0010110000111" => index <= 6;
         when "0010110001000" => index <= 8;
         when "0010110001001" => index <= 7;
         when "0010110001010" => index <= 7;
         when "0010110001011" => index <= 6;
         when "0010110001100" => index <= 7;
         when "0010110001101" => index <= 6;
         when "0010110001110" => index <= 6;
         when "0010110001111" => index <= 5;
         when "0010110010000" => index <= 8;
         when "0010110010001" => index <= 7;
         when "0010110010010" => index <= 7;
         when "0010110010011" => index <= 6;
         when "0010110010100" => index <= 7;
         when "0010110010101" => index <= 6;
         when "0010110010110" => index <= 6;
         when "0010110010111" => index <= 6;
         when "0010110011000" => index <= 7;
         when "0010110011001" => index <= 6;
         when "0010110011010" => index <= 6;
         when "0010110011011" => index <= 6;
         when "0010110011100" => index <= 7;
         when "0010110011101" => index <= 6;
         when "0010110011110" => index <= 6;
         when "0010110011111" => index <= 5;
         when "0010110100000" => index <= 8;
         when "0010110100001" => index <= 7;
         when "0010110100010" => index <= 7;
         when "0010110100011" => index <= 6;
         when "0010110100100" => index <= 7;
         when "0010110100101" => index <= 6;
         when "0010110100110" => index <= 6;
         when "0010110100111" => index <= 6;
         when "0010110101000" => index <= 8;
         when "0010110101001" => index <= 6;
         when "0010110101010" => index <= 7;
         when "0010110101011" => index <= 6;
         when "0010110101100" => index <= 7;
         when "0010110101101" => index <= 6;
         when "0010110101110" => index <= 6;
         when "0010110101111" => index <= 6;
         when "0010110110000" => index <= 8;
         when "0010110110001" => index <= 7;
         when "0010110110010" => index <= 7;
         when "0010110110011" => index <= 6;
         when "0010110110100" => index <= 7;
         when "0010110110101" => index <= 6;
         when "0010110110110" => index <= 6;
         when "0010110110111" => index <= 6;
         when "0010110111000" => index <= 7;
         when "0010110111001" => index <= 6;
         when "0010110111010" => index <= 6;
         when "0010110111011" => index <= 6;
         when "0010110111100" => index <= 7;
         when "0010110111101" => index <= 6;
         when "0010110111110" => index <= 6;
         when "0010110111111" => index <= 5;
         when "0010111000000" => index <= 9;
         when "0010111000001" => index <= 7;
         when "0010111000010" => index <= 7;
         when "0010111000011" => index <= 6;
         when "0010111000100" => index <= 8;
         when "0010111000101" => index <= 6;
         when "0010111000110" => index <= 7;
         when "0010111000111" => index <= 6;
         when "0010111001000" => index <= 8;
         when "0010111001001" => index <= 7;
         when "0010111001010" => index <= 7;
         when "0010111001011" => index <= 6;
         when "0010111001100" => index <= 7;
         when "0010111001101" => index <= 6;
         when "0010111001110" => index <= 6;
         when "0010111001111" => index <= 6;
         when "0010111010000" => index <= 8;
         when "0010111010001" => index <= 7;
         when "0010111010010" => index <= 7;
         when "0010111010011" => index <= 6;
         when "0010111010100" => index <= 7;
         when "0010111010101" => index <= 6;
         when "0010111010110" => index <= 6;
         when "0010111010111" => index <= 6;
         when "0010111011000" => index <= 7;
         when "0010111011001" => index <= 6;
         when "0010111011010" => index <= 7;
         when "0010111011011" => index <= 6;
         when "0010111011100" => index <= 7;
         when "0010111011101" => index <= 6;
         when "0010111011110" => index <= 6;
         when "0010111011111" => index <= 6;
         when "0010111100000" => index <= 8;
         when "0010111100001" => index <= 7;
         when "0010111100010" => index <= 7;
         when "0010111100011" => index <= 6;
         when "0010111100100" => index <= 7;
         when "0010111100101" => index <= 6;
         when "0010111100110" => index <= 7;
         when "0010111100111" => index <= 6;
         when "0010111101000" => index <= 8;
         when "0010111101001" => index <= 7;
         when "0010111101010" => index <= 7;
         when "0010111101011" => index <= 6;
         when "0010111101100" => index <= 7;
         when "0010111101101" => index <= 6;
         when "0010111101110" => index <= 6;
         when "0010111101111" => index <= 6;
         when "0010111110000" => index <= 8;
         when "0010111110001" => index <= 7;
         when "0010111110010" => index <= 7;
         when "0010111110011" => index <= 6;
         when "0010111110100" => index <= 7;
         when "0010111110101" => index <= 6;
         when "0010111110110" => index <= 6;
         when "0010111110111" => index <= 6;
         when "0010111111000" => index <= 7;
         when "0010111111001" => index <= 6;
         when "0010111111010" => index <= 6;
         when "0010111111011" => index <= 6;
         when "0010111111100" => index <= 7;
         when "0010111111101" => index <= 6;
         when "0010111111110" => index <= 6;
         when "0010111111111" => index <= 6;
         when "0011000000000" => index <= 10;
         when "0011000000001" => index <= 7;
         when "0011000000010" => index <= 8;
         when "0011000000011" => index <= 6;
         when "0011000000100" => index <= 8;
         when "0011000000101" => index <= 6;
         when "0011000000110" => index <= 6;
         when "0011000000111" => index <= 5;
         when "0011000001000" => index <= 8;
         when "0011000001001" => index <= 6;
         when "0011000001010" => index <= 7;
         when "0011000001011" => index <= 6;
         when "0011000001100" => index <= 7;
         when "0011000001101" => index <= 6;
         when "0011000001110" => index <= 6;
         when "0011000001111" => index <= 5;
         when "0011000010000" => index <= 9;
         when "0011000010001" => index <= 7;
         when "0011000010010" => index <= 7;
         when "0011000010011" => index <= 6;
         when "0011000010100" => index <= 7;
         when "0011000010101" => index <= 6;
         when "0011000010110" => index <= 6;
         when "0011000010111" => index <= 5;
         when "0011000011000" => index <= 8;
         when "0011000011001" => index <= 6;
         when "0011000011010" => index <= 6;
         when "0011000011011" => index <= 6;
         when "0011000011100" => index <= 7;
         when "0011000011101" => index <= 6;
         when "0011000011110" => index <= 6;
         when "0011000011111" => index <= 5;
         when "0011000100000" => index <= 9;
         when "0011000100001" => index <= 7;
         when "0011000100010" => index <= 7;
         when "0011000100011" => index <= 6;
         when "0011000100100" => index <= 8;
         when "0011000100101" => index <= 6;
         when "0011000100110" => index <= 6;
         when "0011000100111" => index <= 6;
         when "0011000101000" => index <= 8;
         when "0011000101001" => index <= 6;
         when "0011000101010" => index <= 7;
         when "0011000101011" => index <= 6;
         when "0011000101100" => index <= 7;
         when "0011000101101" => index <= 6;
         when "0011000101110" => index <= 6;
         when "0011000101111" => index <= 5;
         when "0011000110000" => index <= 8;
         when "0011000110001" => index <= 7;
         when "0011000110010" => index <= 7;
         when "0011000110011" => index <= 6;
         when "0011000110100" => index <= 7;
         when "0011000110101" => index <= 6;
         when "0011000110110" => index <= 6;
         when "0011000110111" => index <= 5;
         when "0011000111000" => index <= 7;
         when "0011000111001" => index <= 6;
         when "0011000111010" => index <= 6;
         when "0011000111011" => index <= 6;
         when "0011000111100" => index <= 6;
         when "0011000111101" => index <= 6;
         when "0011000111110" => index <= 6;
         when "0011000111111" => index <= 5;
         when "0011001000000" => index <= 9;
         when "0011001000001" => index <= 7;
         when "0011001000010" => index <= 8;
         when "0011001000011" => index <= 6;
         when "0011001000100" => index <= 8;
         when "0011001000101" => index <= 6;
         when "0011001000110" => index <= 7;
         when "0011001000111" => index <= 6;
         when "0011001001000" => index <= 8;
         when "0011001001001" => index <= 7;
         when "0011001001010" => index <= 7;
         when "0011001001011" => index <= 6;
         when "0011001001100" => index <= 7;
         when "0011001001101" => index <= 6;
         when "0011001001110" => index <= 6;
         when "0011001001111" => index <= 5;
         when "0011001010000" => index <= 8;
         when "0011001010001" => index <= 7;
         when "0011001010010" => index <= 7;
         when "0011001010011" => index <= 6;
         when "0011001010100" => index <= 7;
         when "0011001010101" => index <= 6;
         when "0011001010110" => index <= 6;
         when "0011001010111" => index <= 6;
         when "0011001011000" => index <= 7;
         when "0011001011001" => index <= 6;
         when "0011001011010" => index <= 6;
         when "0011001011011" => index <= 6;
         when "0011001011100" => index <= 7;
         when "0011001011101" => index <= 6;
         when "0011001011110" => index <= 6;
         when "0011001011111" => index <= 5;
         when "0011001100000" => index <= 8;
         when "0011001100001" => index <= 7;
         when "0011001100010" => index <= 7;
         when "0011001100011" => index <= 6;
         when "0011001100100" => index <= 7;
         when "0011001100101" => index <= 6;
         when "0011001100110" => index <= 6;
         when "0011001100111" => index <= 6;
         when "0011001101000" => index <= 8;
         when "0011001101001" => index <= 6;
         when "0011001101010" => index <= 7;
         when "0011001101011" => index <= 6;
         when "0011001101100" => index <= 7;
         when "0011001101101" => index <= 6;
         when "0011001101110" => index <= 6;
         when "0011001101111" => index <= 6;
         when "0011001110000" => index <= 8;
         when "0011001110001" => index <= 7;
         when "0011001110010" => index <= 7;
         when "0011001110011" => index <= 6;
         when "0011001110100" => index <= 7;
         when "0011001110101" => index <= 6;
         when "0011001110110" => index <= 6;
         when "0011001110111" => index <= 6;
         when "0011001111000" => index <= 7;
         when "0011001111001" => index <= 6;
         when "0011001111010" => index <= 6;
         when "0011001111011" => index <= 6;
         when "0011001111100" => index <= 7;
         when "0011001111101" => index <= 6;
         when "0011001111110" => index <= 6;
         when "0011001111111" => index <= 5;
         when "0011010000000" => index <= 10;
         when "0011010000001" => index <= 8;
         when "0011010000010" => index <= 8;
         when "0011010000011" => index <= 6;
         when "0011010000100" => index <= 8;
         when "0011010000101" => index <= 7;
         when "0011010000110" => index <= 7;
         when "0011010000111" => index <= 6;
         when "0011010001000" => index <= 8;
         when "0011010001001" => index <= 7;
         when "0011010001010" => index <= 7;
         when "0011010001011" => index <= 6;
         when "0011010001100" => index <= 7;
         when "0011010001101" => index <= 6;
         when "0011010001110" => index <= 6;
         when "0011010001111" => index <= 6;
         when "0011010010000" => index <= 8;
         when "0011010010001" => index <= 7;
         when "0011010010010" => index <= 7;
         when "0011010010011" => index <= 6;
         when "0011010010100" => index <= 7;
         when "0011010010101" => index <= 6;
         when "0011010010110" => index <= 6;
         when "0011010010111" => index <= 6;
         when "0011010011000" => index <= 8;
         when "0011010011001" => index <= 6;
         when "0011010011010" => index <= 7;
         when "0011010011011" => index <= 6;
         when "0011010011100" => index <= 7;
         when "0011010011101" => index <= 6;
         when "0011010011110" => index <= 6;
         when "0011010011111" => index <= 6;
         when "0011010100000" => index <= 9;
         when "0011010100001" => index <= 7;
         when "0011010100010" => index <= 7;
         when "0011010100011" => index <= 6;
         when "0011010100100" => index <= 8;
         when "0011010100101" => index <= 6;
         when "0011010100110" => index <= 7;
         when "0011010100111" => index <= 6;
         when "0011010101000" => index <= 8;
         when "0011010101001" => index <= 7;
         when "0011010101010" => index <= 7;
         when "0011010101011" => index <= 6;
         when "0011010101100" => index <= 7;
         when "0011010101101" => index <= 6;
         when "0011010101110" => index <= 6;
         when "0011010101111" => index <= 6;
         when "0011010110000" => index <= 8;
         when "0011010110001" => index <= 7;
         when "0011010110010" => index <= 7;
         when "0011010110011" => index <= 6;
         when "0011010110100" => index <= 7;
         when "0011010110101" => index <= 6;
         when "0011010110110" => index <= 6;
         when "0011010110111" => index <= 6;
         when "0011010111000" => index <= 7;
         when "0011010111001" => index <= 6;
         when "0011010111010" => index <= 7;
         when "0011010111011" => index <= 6;
         when "0011010111100" => index <= 7;
         when "0011010111101" => index <= 6;
         when "0011010111110" => index <= 6;
         when "0011010111111" => index <= 6;
         when "0011011000000" => index <= 9;
         when "0011011000001" => index <= 7;
         when "0011011000010" => index <= 8;
         when "0011011000011" => index <= 6;
         when "0011011000100" => index <= 8;
         when "0011011000101" => index <= 7;
         when "0011011000110" => index <= 7;
         when "0011011000111" => index <= 6;
         when "0011011001000" => index <= 8;
         when "0011011001001" => index <= 7;
         when "0011011001010" => index <= 7;
         when "0011011001011" => index <= 6;
         when "0011011001100" => index <= 7;
         when "0011011001101" => index <= 6;
         when "0011011001110" => index <= 6;
         when "0011011001111" => index <= 6;
         when "0011011010000" => index <= 8;
         when "0011011010001" => index <= 7;
         when "0011011010010" => index <= 7;
         when "0011011010011" => index <= 6;
         when "0011011010100" => index <= 7;
         when "0011011010101" => index <= 6;
         when "0011011010110" => index <= 7;
         when "0011011010111" => index <= 6;
         when "0011011011000" => index <= 8;
         when "0011011011001" => index <= 7;
         when "0011011011010" => index <= 7;
         when "0011011011011" => index <= 6;
         when "0011011011100" => index <= 7;
         when "0011011011101" => index <= 6;
         when "0011011011110" => index <= 6;
         when "0011011011111" => index <= 6;
         when "0011011100000" => index <= 8;
         when "0011011100001" => index <= 7;
         when "0011011100010" => index <= 7;
         when "0011011100011" => index <= 6;
         when "0011011100100" => index <= 8;
         when "0011011100101" => index <= 7;
         when "0011011100110" => index <= 7;
         when "0011011100111" => index <= 6;
         when "0011011101000" => index <= 8;
         when "0011011101001" => index <= 7;
         when "0011011101010" => index <= 7;
         when "0011011101011" => index <= 6;
         when "0011011101100" => index <= 7;
         when "0011011101101" => index <= 6;
         when "0011011101110" => index <= 6;
         when "0011011101111" => index <= 6;
         when "0011011110000" => index <= 8;
         when "0011011110001" => index <= 7;
         when "0011011110010" => index <= 7;
         when "0011011110011" => index <= 6;
         when "0011011110100" => index <= 7;
         when "0011011110101" => index <= 6;
         when "0011011110110" => index <= 6;
         when "0011011110111" => index <= 6;
         when "0011011111000" => index <= 7;
         when "0011011111001" => index <= 6;
         when "0011011111010" => index <= 7;
         when "0011011111011" => index <= 6;
         when "0011011111100" => index <= 7;
         when "0011011111101" => index <= 6;
         when "0011011111110" => index <= 6;
         when "0011011111111" => index <= 6;
         when "0011100000000" => index <= 10;
         when "0011100000001" => index <= 8;
         when "0011100000010" => index <= 8;
         when "0011100000011" => index <= 7;
         when "0011100000100" => index <= 8;
         when "0011100000101" => index <= 7;
         when "0011100000110" => index <= 7;
         when "0011100000111" => index <= 6;
         when "0011100001000" => index <= 8;
         when "0011100001001" => index <= 7;
         when "0011100001010" => index <= 7;
         when "0011100001011" => index <= 6;
         when "0011100001100" => index <= 7;
         when "0011100001101" => index <= 6;
         when "0011100001110" => index <= 6;
         when "0011100001111" => index <= 6;
         when "0011100010000" => index <= 9;
         when "0011100010001" => index <= 7;
         when "0011100010010" => index <= 7;
         when "0011100010011" => index <= 6;
         when "0011100010100" => index <= 8;
         when "0011100010101" => index <= 6;
         when "0011100010110" => index <= 7;
         when "0011100010111" => index <= 6;
         when "0011100011000" => index <= 8;
         when "0011100011001" => index <= 7;
         when "0011100011010" => index <= 7;
         when "0011100011011" => index <= 6;
         when "0011100011100" => index <= 7;
         when "0011100011101" => index <= 6;
         when "0011100011110" => index <= 6;
         when "0011100011111" => index <= 6;
         when "0011100100000" => index <= 9;
         when "0011100100001" => index <= 7;
         when "0011100100010" => index <= 8;
         when "0011100100011" => index <= 6;
         when "0011100100100" => index <= 8;
         when "0011100100101" => index <= 7;
         when "0011100100110" => index <= 7;
         when "0011100100111" => index <= 6;
         when "0011100101000" => index <= 8;
         when "0011100101001" => index <= 7;
         when "0011100101010" => index <= 7;
         when "0011100101011" => index <= 6;
         when "0011100101100" => index <= 7;
         when "0011100101101" => index <= 6;
         when "0011100101110" => index <= 6;
         when "0011100101111" => index <= 6;
         when "0011100110000" => index <= 8;
         when "0011100110001" => index <= 7;
         when "0011100110010" => index <= 7;
         when "0011100110011" => index <= 6;
         when "0011100110100" => index <= 7;
         when "0011100110101" => index <= 6;
         when "0011100110110" => index <= 7;
         when "0011100110111" => index <= 6;
         when "0011100111000" => index <= 8;
         when "0011100111001" => index <= 7;
         when "0011100111010" => index <= 7;
         when "0011100111011" => index <= 6;
         when "0011100111100" => index <= 7;
         when "0011100111101" => index <= 6;
         when "0011100111110" => index <= 6;
         when "0011100111111" => index <= 6;
         when "0011101000000" => index <= 9;
         when "0011101000001" => index <= 8;
         when "0011101000010" => index <= 8;
         when "0011101000011" => index <= 7;
         when "0011101000100" => index <= 8;
         when "0011101000101" => index <= 7;
         when "0011101000110" => index <= 7;
         when "0011101000111" => index <= 6;
         when "0011101001000" => index <= 8;
         when "0011101001001" => index <= 7;
         when "0011101001010" => index <= 7;
         when "0011101001011" => index <= 6;
         when "0011101001100" => index <= 7;
         when "0011101001101" => index <= 6;
         when "0011101001110" => index <= 7;
         when "0011101001111" => index <= 6;
         when "0011101010000" => index <= 8;
         when "0011101010001" => index <= 7;
         when "0011101010010" => index <= 7;
         when "0011101010011" => index <= 6;
         when "0011101010100" => index <= 8;
         when "0011101010101" => index <= 7;
         when "0011101010110" => index <= 7;
         when "0011101010111" => index <= 6;
         when "0011101011000" => index <= 8;
         when "0011101011001" => index <= 7;
         when "0011101011010" => index <= 7;
         when "0011101011011" => index <= 6;
         when "0011101011100" => index <= 7;
         when "0011101011101" => index <= 6;
         when "0011101011110" => index <= 6;
         when "0011101011111" => index <= 6;
         when "0011101100000" => index <= 9;
         when "0011101100001" => index <= 7;
         when "0011101100010" => index <= 8;
         when "0011101100011" => index <= 7;
         when "0011101100100" => index <= 8;
         when "0011101100101" => index <= 7;
         when "0011101100110" => index <= 7;
         when "0011101100111" => index <= 6;
         when "0011101101000" => index <= 8;
         when "0011101101001" => index <= 7;
         when "0011101101010" => index <= 7;
         when "0011101101011" => index <= 6;
         when "0011101101100" => index <= 7;
         when "0011101101101" => index <= 6;
         when "0011101101110" => index <= 6;
         when "0011101101111" => index <= 6;
         when "0011101110000" => index <= 8;
         when "0011101110001" => index <= 7;
         when "0011101110010" => index <= 7;
         when "0011101110011" => index <= 6;
         when "0011101110100" => index <= 7;
         when "0011101110101" => index <= 6;
         when "0011101110110" => index <= 7;
         when "0011101110111" => index <= 6;
         when "0011101111000" => index <= 7;
         when "0011101111001" => index <= 7;
         when "0011101111010" => index <= 7;
         when "0011101111011" => index <= 6;
         when "0011101111100" => index <= 7;
         when "0011101111101" => index <= 6;
         when "0011101111110" => index <= 6;
         when "0011101111111" => index <= 6;
         when "0011110000000" => index <= 10;
         when "0011110000001" => index <= 8;
         when "0011110000010" => index <= 8;
         when "0011110000011" => index <= 7;
         when "0011110000100" => index <= 8;
         when "0011110000101" => index <= 7;
         when "0011110000110" => index <= 7;
         when "0011110000111" => index <= 6;
         when "0011110001000" => index <= 8;
         when "0011110001001" => index <= 7;
         when "0011110001010" => index <= 7;
         when "0011110001011" => index <= 6;
         when "0011110001100" => index <= 8;
         when "0011110001101" => index <= 7;
         when "0011110001110" => index <= 7;
         when "0011110001111" => index <= 6;
         when "0011110010000" => index <= 9;
         when "0011110010001" => index <= 7;
         when "0011110010010" => index <= 8;
         when "0011110010011" => index <= 7;
         when "0011110010100" => index <= 8;
         when "0011110010101" => index <= 7;
         when "0011110010110" => index <= 7;
         when "0011110010111" => index <= 6;
         when "0011110011000" => index <= 8;
         when "0011110011001" => index <= 7;
         when "0011110011010" => index <= 7;
         when "0011110011011" => index <= 6;
         when "0011110011100" => index <= 7;
         when "0011110011101" => index <= 6;
         when "0011110011110" => index <= 6;
         when "0011110011111" => index <= 6;
         when "0011110100000" => index <= 9;
         when "0011110100001" => index <= 8;
         when "0011110100010" => index <= 8;
         when "0011110100011" => index <= 7;
         when "0011110100100" => index <= 8;
         when "0011110100101" => index <= 7;
         when "0011110100110" => index <= 7;
         when "0011110100111" => index <= 6;
         when "0011110101000" => index <= 8;
         when "0011110101001" => index <= 7;
         when "0011110101010" => index <= 7;
         when "0011110101011" => index <= 6;
         when "0011110101100" => index <= 7;
         when "0011110101101" => index <= 6;
         when "0011110101110" => index <= 7;
         when "0011110101111" => index <= 6;
         when "0011110110000" => index <= 8;
         when "0011110110001" => index <= 7;
         when "0011110110010" => index <= 7;
         when "0011110110011" => index <= 6;
         when "0011110110100" => index <= 7;
         when "0011110110101" => index <= 7;
         when "0011110110110" => index <= 7;
         when "0011110110111" => index <= 6;
         when "0011110111000" => index <= 8;
         when "0011110111001" => index <= 7;
         when "0011110111010" => index <= 7;
         when "0011110111011" => index <= 6;
         when "0011110111100" => index <= 7;
         when "0011110111101" => index <= 6;
         when "0011110111110" => index <= 6;
         when "0011110111111" => index <= 6;
         when "0011111000000" => index <= 9;
         when "0011111000001" => index <= 8;
         when "0011111000010" => index <= 8;
         when "0011111000011" => index <= 7;
         when "0011111000100" => index <= 8;
         when "0011111000101" => index <= 7;
         when "0011111000110" => index <= 7;
         when "0011111000111" => index <= 6;
         when "0011111001000" => index <= 8;
         when "0011111001001" => index <= 7;
         when "0011111001010" => index <= 7;
         when "0011111001011" => index <= 6;
         when "0011111001100" => index <= 7;
         when "0011111001101" => index <= 7;
         when "0011111001110" => index <= 7;
         when "0011111001111" => index <= 6;
         when "0011111010000" => index <= 8;
         when "0011111010001" => index <= 7;
         when "0011111010010" => index <= 7;
         when "0011111010011" => index <= 7;
         when "0011111010100" => index <= 8;
         when "0011111010101" => index <= 7;
         when "0011111010110" => index <= 7;
         when "0011111010111" => index <= 6;
         when "0011111011000" => index <= 8;
         when "0011111011001" => index <= 7;
         when "0011111011010" => index <= 7;
         when "0011111011011" => index <= 6;
         when "0011111011100" => index <= 7;
         when "0011111011101" => index <= 6;
         when "0011111011110" => index <= 7;
         when "0011111011111" => index <= 6;
         when "0011111100000" => index <= 8;
         when "0011111100001" => index <= 7;
         when "0011111100010" => index <= 8;
         when "0011111100011" => index <= 7;
         when "0011111100100" => index <= 8;
         when "0011111100101" => index <= 7;
         when "0011111100110" => index <= 7;
         when "0011111100111" => index <= 6;
         when "0011111101000" => index <= 8;
         when "0011111101001" => index <= 7;
         when "0011111101010" => index <= 7;
         when "0011111101011" => index <= 6;
         when "0011111101100" => index <= 7;
         when "0011111101101" => index <= 7;
         when "0011111101110" => index <= 7;
         when "0011111101111" => index <= 6;
         when "0011111110000" => index <= 8;
         when "0011111110001" => index <= 7;
         when "0011111110010" => index <= 7;
         when "0011111110011" => index <= 7;
         when "0011111110100" => index <= 7;
         when "0011111110101" => index <= 7;
         when "0011111110110" => index <= 7;
         when "0011111110111" => index <= 6;
         when "0011111111000" => index <= 8;
         when "0011111111001" => index <= 7;
         when "0011111111010" => index <= 7;
         when "0011111111011" => index <= 6;
         when "0011111111100" => index <= 7;
         when "0011111111101" => index <= 6;
         when "0011111111110" => index <= 6;
         when "0011111111111" => index <= 6;
         when "0100000000000" => index <= 12;
         when "0100000000001" => index <= 6;
         when "0100000000010" => index <= 7;
         when "0100000000011" => index <= 5;
         when "0100000000100" => index <= 8;
         when "0100000000101" => index <= 5;
         when "0100000000110" => index <= 6;
         when "0100000000111" => index <= 4;
         when "0100000001000" => index <= 8;
         when "0100000001001" => index <= 6;
         when "0100000001010" => index <= 6;
         when "0100000001011" => index <= 5;
         when "0100000001100" => index <= 6;
         when "0100000001101" => index <= 5;
         when "0100000001110" => index <= 5;
         when "0100000001111" => index <= 4;
         when "0100000010000" => index <= 8;
         when "0100000010001" => index <= 6;
         when "0100000010010" => index <= 6;
         when "0100000010011" => index <= 5;
         when "0100000010100" => index <= 7;
         when "0100000010101" => index <= 5;
         when "0100000010110" => index <= 6;
         when "0100000010111" => index <= 5;
         when "0100000011000" => index <= 7;
         when "0100000011001" => index <= 6;
         when "0100000011010" => index <= 6;
         when "0100000011011" => index <= 5;
         when "0100000011100" => index <= 6;
         when "0100000011101" => index <= 5;
         when "0100000011110" => index <= 5;
         when "0100000011111" => index <= 4;
         when "0100000100000" => index <= 9;
         when "0100000100001" => index <= 6;
         when "0100000100010" => index <= 7;
         when "0100000100011" => index <= 5;
         when "0100000100100" => index <= 7;
         when "0100000100101" => index <= 6;
         when "0100000100110" => index <= 6;
         when "0100000100111" => index <= 5;
         when "0100000101000" => index <= 7;
         when "0100000101001" => index <= 6;
         when "0100000101010" => index <= 6;
         when "0100000101011" => index <= 5;
         when "0100000101100" => index <= 6;
         when "0100000101101" => index <= 5;
         when "0100000101110" => index <= 5;
         when "0100000101111" => index <= 5;
         when "0100000110000" => index <= 8;
         when "0100000110001" => index <= 6;
         when "0100000110010" => index <= 6;
         when "0100000110011" => index <= 5;
         when "0100000110100" => index <= 6;
         when "0100000110101" => index <= 5;
         when "0100000110110" => index <= 6;
         when "0100000110111" => index <= 5;
         when "0100000111000" => index <= 7;
         when "0100000111001" => index <= 6;
         when "0100000111010" => index <= 6;
         when "0100000111011" => index <= 5;
         when "0100000111100" => index <= 6;
         when "0100000111101" => index <= 5;
         when "0100000111110" => index <= 5;
         when "0100000111111" => index <= 5;
         when "0100001000000" => index <= 10;
         when "0100001000001" => index <= 7;
         when "0100001000010" => index <= 7;
         when "0100001000011" => index <= 6;
         when "0100001000100" => index <= 7;
         when "0100001000101" => index <= 6;
         when "0100001000110" => index <= 6;
         when "0100001000111" => index <= 5;
         when "0100001001000" => index <= 8;
         when "0100001001001" => index <= 6;
         when "0100001001010" => index <= 6;
         when "0100001001011" => index <= 5;
         when "0100001001100" => index <= 6;
         when "0100001001101" => index <= 5;
         when "0100001001110" => index <= 6;
         when "0100001001111" => index <= 5;
         when "0100001010000" => index <= 8;
         when "0100001010001" => index <= 6;
         when "0100001010010" => index <= 6;
         when "0100001010011" => index <= 5;
         when "0100001010100" => index <= 7;
         when "0100001010101" => index <= 6;
         when "0100001010110" => index <= 6;
         when "0100001010111" => index <= 5;
         when "0100001011000" => index <= 7;
         when "0100001011001" => index <= 6;
         when "0100001011010" => index <= 6;
         when "0100001011011" => index <= 5;
         when "0100001011100" => index <= 6;
         when "0100001011101" => index <= 5;
         when "0100001011110" => index <= 6;
         when "0100001011111" => index <= 5;
         when "0100001100000" => index <= 8;
         when "0100001100001" => index <= 6;
         when "0100001100010" => index <= 7;
         when "0100001100011" => index <= 6;
         when "0100001100100" => index <= 7;
         when "0100001100101" => index <= 6;
         when "0100001100110" => index <= 6;
         when "0100001100111" => index <= 5;
         when "0100001101000" => index <= 7;
         when "0100001101001" => index <= 6;
         when "0100001101010" => index <= 6;
         when "0100001101011" => index <= 5;
         when "0100001101100" => index <= 6;
         when "0100001101101" => index <= 6;
         when "0100001101110" => index <= 6;
         when "0100001101111" => index <= 5;
         when "0100001110000" => index <= 8;
         when "0100001110001" => index <= 6;
         when "0100001110010" => index <= 6;
         when "0100001110011" => index <= 6;
         when "0100001110100" => index <= 7;
         when "0100001110101" => index <= 6;
         when "0100001110110" => index <= 6;
         when "0100001110111" => index <= 5;
         when "0100001111000" => index <= 7;
         when "0100001111001" => index <= 6;
         when "0100001111010" => index <= 6;
         when "0100001111011" => index <= 5;
         when "0100001111100" => index <= 6;
         when "0100001111101" => index <= 5;
         when "0100001111110" => index <= 6;
         when "0100001111111" => index <= 5;
         when "0100010000000" => index <= 10;
         when "0100010000001" => index <= 7;
         when "0100010000010" => index <= 7;
         when "0100010000011" => index <= 6;
         when "0100010000100" => index <= 8;
         when "0100010000101" => index <= 6;
         when "0100010000110" => index <= 6;
         when "0100010000111" => index <= 5;
         when "0100010001000" => index <= 8;
         when "0100010001001" => index <= 6;
         when "0100010001010" => index <= 6;
         when "0100010001011" => index <= 5;
         when "0100010001100" => index <= 7;
         when "0100010001101" => index <= 6;
         when "0100010001110" => index <= 6;
         when "0100010001111" => index <= 5;
         when "0100010010000" => index <= 8;
         when "0100010010001" => index <= 6;
         when "0100010010010" => index <= 7;
         when "0100010010011" => index <= 6;
         when "0100010010100" => index <= 7;
         when "0100010010101" => index <= 6;
         when "0100010010110" => index <= 6;
         when "0100010010111" => index <= 5;
         when "0100010011000" => index <= 7;
         when "0100010011001" => index <= 6;
         when "0100010011010" => index <= 6;
         when "0100010011011" => index <= 5;
         when "0100010011100" => index <= 6;
         when "0100010011101" => index <= 6;
         when "0100010011110" => index <= 6;
         when "0100010011111" => index <= 5;
         when "0100010100000" => index <= 9;
         when "0100010100001" => index <= 7;
         when "0100010100010" => index <= 7;
         when "0100010100011" => index <= 6;
         when "0100010100100" => index <= 7;
         when "0100010100101" => index <= 6;
         when "0100010100110" => index <= 6;
         when "0100010100111" => index <= 5;
         when "0100010101000" => index <= 8;
         when "0100010101001" => index <= 6;
         when "0100010101010" => index <= 6;
         when "0100010101011" => index <= 6;
         when "0100010101100" => index <= 7;
         when "0100010101101" => index <= 6;
         when "0100010101110" => index <= 6;
         when "0100010101111" => index <= 5;
         when "0100010110000" => index <= 8;
         when "0100010110001" => index <= 6;
         when "0100010110010" => index <= 7;
         when "0100010110011" => index <= 6;
         when "0100010110100" => index <= 7;
         when "0100010110101" => index <= 6;
         when "0100010110110" => index <= 6;
         when "0100010110111" => index <= 5;
         when "0100010111000" => index <= 7;
         when "0100010111001" => index <= 6;
         when "0100010111010" => index <= 6;
         when "0100010111011" => index <= 5;
         when "0100010111100" => index <= 6;
         when "0100010111101" => index <= 6;
         when "0100010111110" => index <= 6;
         when "0100010111111" => index <= 5;
         when "0100011000000" => index <= 9;
         when "0100011000001" => index <= 7;
         when "0100011000010" => index <= 7;
         when "0100011000011" => index <= 6;
         when "0100011000100" => index <= 8;
         when "0100011000101" => index <= 6;
         when "0100011000110" => index <= 6;
         when "0100011000111" => index <= 6;
         when "0100011001000" => index <= 8;
         when "0100011001001" => index <= 6;
         when "0100011001010" => index <= 7;
         when "0100011001011" => index <= 6;
         when "0100011001100" => index <= 7;
         when "0100011001101" => index <= 6;
         when "0100011001110" => index <= 6;
         when "0100011001111" => index <= 5;
         when "0100011010000" => index <= 8;
         when "0100011010001" => index <= 7;
         when "0100011010010" => index <= 7;
         when "0100011010011" => index <= 6;
         when "0100011010100" => index <= 7;
         when "0100011010101" => index <= 6;
         when "0100011010110" => index <= 6;
         when "0100011010111" => index <= 5;
         when "0100011011000" => index <= 7;
         when "0100011011001" => index <= 6;
         when "0100011011010" => index <= 6;
         when "0100011011011" => index <= 6;
         when "0100011011100" => index <= 6;
         when "0100011011101" => index <= 6;
         when "0100011011110" => index <= 6;
         when "0100011011111" => index <= 5;
         when "0100011100000" => index <= 8;
         when "0100011100001" => index <= 7;
         when "0100011100010" => index <= 7;
         when "0100011100011" => index <= 6;
         when "0100011100100" => index <= 7;
         when "0100011100101" => index <= 6;
         when "0100011100110" => index <= 6;
         when "0100011100111" => index <= 6;
         when "0100011101000" => index <= 7;
         when "0100011101001" => index <= 6;
         when "0100011101010" => index <= 6;
         when "0100011101011" => index <= 6;
         when "0100011101100" => index <= 7;
         when "0100011101101" => index <= 6;
         when "0100011101110" => index <= 6;
         when "0100011101111" => index <= 5;
         when "0100011110000" => index <= 8;
         when "0100011110001" => index <= 6;
         when "0100011110010" => index <= 7;
         when "0100011110011" => index <= 6;
         when "0100011110100" => index <= 7;
         when "0100011110101" => index <= 6;
         when "0100011110110" => index <= 6;
         when "0100011110111" => index <= 6;
         when "0100011111000" => index <= 7;
         when "0100011111001" => index <= 6;
         when "0100011111010" => index <= 6;
         when "0100011111011" => index <= 6;
         when "0100011111100" => index <= 6;
         when "0100011111101" => index <= 6;
         when "0100011111110" => index <= 6;
         when "0100011111111" => index <= 5;
         when "0100100000000" => index <= 10;
         when "0100100000001" => index <= 7;
         when "0100100000010" => index <= 8;
         when "0100100000011" => index <= 6;
         when "0100100000100" => index <= 8;
         when "0100100000101" => index <= 6;
         when "0100100000110" => index <= 6;
         when "0100100000111" => index <= 5;
         when "0100100001000" => index <= 8;
         when "0100100001001" => index <= 6;
         when "0100100001010" => index <= 7;
         when "0100100001011" => index <= 6;
         when "0100100001100" => index <= 7;
         when "0100100001101" => index <= 6;
         when "0100100001110" => index <= 6;
         when "0100100001111" => index <= 5;
         when "0100100010000" => index <= 9;
         when "0100100010001" => index <= 7;
         when "0100100010010" => index <= 7;
         when "0100100010011" => index <= 6;
         when "0100100010100" => index <= 7;
         when "0100100010101" => index <= 6;
         when "0100100010110" => index <= 6;
         when "0100100010111" => index <= 5;
         when "0100100011000" => index <= 8;
         when "0100100011001" => index <= 6;
         when "0100100011010" => index <= 6;
         when "0100100011011" => index <= 6;
         when "0100100011100" => index <= 7;
         when "0100100011101" => index <= 6;
         when "0100100011110" => index <= 6;
         when "0100100011111" => index <= 5;
         when "0100100100000" => index <= 9;
         when "0100100100001" => index <= 7;
         when "0100100100010" => index <= 7;
         when "0100100100011" => index <= 6;
         when "0100100100100" => index <= 8;
         when "0100100100101" => index <= 6;
         when "0100100100110" => index <= 6;
         when "0100100100111" => index <= 6;
         when "0100100101000" => index <= 8;
         when "0100100101001" => index <= 6;
         when "0100100101010" => index <= 7;
         when "0100100101011" => index <= 6;
         when "0100100101100" => index <= 7;
         when "0100100101101" => index <= 6;
         when "0100100101110" => index <= 6;
         when "0100100101111" => index <= 5;
         when "0100100110000" => index <= 8;
         when "0100100110001" => index <= 7;
         when "0100100110010" => index <= 7;
         when "0100100110011" => index <= 6;
         when "0100100110100" => index <= 7;
         when "0100100110101" => index <= 6;
         when "0100100110110" => index <= 6;
         when "0100100110111" => index <= 5;
         when "0100100111000" => index <= 7;
         when "0100100111001" => index <= 6;
         when "0100100111010" => index <= 6;
         when "0100100111011" => index <= 6;
         when "0100100111100" => index <= 6;
         when "0100100111101" => index <= 6;
         when "0100100111110" => index <= 6;
         when "0100100111111" => index <= 5;
         when "0100101000000" => index <= 9;
         when "0100101000001" => index <= 7;
         when "0100101000010" => index <= 8;
         when "0100101000011" => index <= 6;
         when "0100101000100" => index <= 8;
         when "0100101000101" => index <= 6;
         when "0100101000110" => index <= 7;
         when "0100101000111" => index <= 6;
         when "0100101001000" => index <= 8;
         when "0100101001001" => index <= 7;
         when "0100101001010" => index <= 7;
         when "0100101001011" => index <= 6;
         when "0100101001100" => index <= 7;
         when "0100101001101" => index <= 6;
         when "0100101001110" => index <= 6;
         when "0100101001111" => index <= 5;
         when "0100101010000" => index <= 8;
         when "0100101010001" => index <= 7;
         when "0100101010010" => index <= 7;
         when "0100101010011" => index <= 6;
         when "0100101010100" => index <= 7;
         when "0100101010101" => index <= 6;
         when "0100101010110" => index <= 6;
         when "0100101010111" => index <= 6;
         when "0100101011000" => index <= 7;
         when "0100101011001" => index <= 6;
         when "0100101011010" => index <= 6;
         when "0100101011011" => index <= 6;
         when "0100101011100" => index <= 7;
         when "0100101011101" => index <= 6;
         when "0100101011110" => index <= 6;
         when "0100101011111" => index <= 5;
         when "0100101100000" => index <= 8;
         when "0100101100001" => index <= 7;
         when "0100101100010" => index <= 7;
         when "0100101100011" => index <= 6;
         when "0100101100100" => index <= 7;
         when "0100101100101" => index <= 6;
         when "0100101100110" => index <= 6;
         when "0100101100111" => index <= 6;
         when "0100101101000" => index <= 8;
         when "0100101101001" => index <= 6;
         when "0100101101010" => index <= 7;
         when "0100101101011" => index <= 6;
         when "0100101101100" => index <= 7;
         when "0100101101101" => index <= 6;
         when "0100101101110" => index <= 6;
         when "0100101101111" => index <= 6;
         when "0100101110000" => index <= 8;
         when "0100101110001" => index <= 7;
         when "0100101110010" => index <= 7;
         when "0100101110011" => index <= 6;
         when "0100101110100" => index <= 7;
         when "0100101110101" => index <= 6;
         when "0100101110110" => index <= 6;
         when "0100101110111" => index <= 6;
         when "0100101111000" => index <= 7;
         when "0100101111001" => index <= 6;
         when "0100101111010" => index <= 6;
         when "0100101111011" => index <= 6;
         when "0100101111100" => index <= 7;
         when "0100101111101" => index <= 6;
         when "0100101111110" => index <= 6;
         when "0100101111111" => index <= 5;
         when "0100110000000" => index <= 10;
         when "0100110000001" => index <= 8;
         when "0100110000010" => index <= 8;
         when "0100110000011" => index <= 6;
         when "0100110000100" => index <= 8;
         when "0100110000101" => index <= 7;
         when "0100110000110" => index <= 7;
         when "0100110000111" => index <= 6;
         when "0100110001000" => index <= 8;
         when "0100110001001" => index <= 7;
         when "0100110001010" => index <= 7;
         when "0100110001011" => index <= 6;
         when "0100110001100" => index <= 7;
         when "0100110001101" => index <= 6;
         when "0100110001110" => index <= 6;
         when "0100110001111" => index <= 6;
         when "0100110010000" => index <= 8;
         when "0100110010001" => index <= 7;
         when "0100110010010" => index <= 7;
         when "0100110010011" => index <= 6;
         when "0100110010100" => index <= 7;
         when "0100110010101" => index <= 6;
         when "0100110010110" => index <= 6;
         when "0100110010111" => index <= 6;
         when "0100110011000" => index <= 8;
         when "0100110011001" => index <= 6;
         when "0100110011010" => index <= 7;
         when "0100110011011" => index <= 6;
         when "0100110011100" => index <= 7;
         when "0100110011101" => index <= 6;
         when "0100110011110" => index <= 6;
         when "0100110011111" => index <= 6;
         when "0100110100000" => index <= 9;
         when "0100110100001" => index <= 7;
         when "0100110100010" => index <= 7;
         when "0100110100011" => index <= 6;
         when "0100110100100" => index <= 8;
         when "0100110100101" => index <= 6;
         when "0100110100110" => index <= 7;
         when "0100110100111" => index <= 6;
         when "0100110101000" => index <= 8;
         when "0100110101001" => index <= 7;
         when "0100110101010" => index <= 7;
         when "0100110101011" => index <= 6;
         when "0100110101100" => index <= 7;
         when "0100110101101" => index <= 6;
         when "0100110101110" => index <= 6;
         when "0100110101111" => index <= 6;
         when "0100110110000" => index <= 8;
         when "0100110110001" => index <= 7;
         when "0100110110010" => index <= 7;
         when "0100110110011" => index <= 6;
         when "0100110110100" => index <= 7;
         when "0100110110101" => index <= 6;
         when "0100110110110" => index <= 6;
         when "0100110110111" => index <= 6;
         when "0100110111000" => index <= 7;
         when "0100110111001" => index <= 6;
         when "0100110111010" => index <= 7;
         when "0100110111011" => index <= 6;
         when "0100110111100" => index <= 7;
         when "0100110111101" => index <= 6;
         when "0100110111110" => index <= 6;
         when "0100110111111" => index <= 6;
         when "0100111000000" => index <= 9;
         when "0100111000001" => index <= 7;
         when "0100111000010" => index <= 8;
         when "0100111000011" => index <= 6;
         when "0100111000100" => index <= 8;
         when "0100111000101" => index <= 7;
         when "0100111000110" => index <= 7;
         when "0100111000111" => index <= 6;
         when "0100111001000" => index <= 8;
         when "0100111001001" => index <= 7;
         when "0100111001010" => index <= 7;
         when "0100111001011" => index <= 6;
         when "0100111001100" => index <= 7;
         when "0100111001101" => index <= 6;
         when "0100111001110" => index <= 6;
         when "0100111001111" => index <= 6;
         when "0100111010000" => index <= 8;
         when "0100111010001" => index <= 7;
         when "0100111010010" => index <= 7;
         when "0100111010011" => index <= 6;
         when "0100111010100" => index <= 7;
         when "0100111010101" => index <= 6;
         when "0100111010110" => index <= 7;
         when "0100111010111" => index <= 6;
         when "0100111011000" => index <= 8;
         when "0100111011001" => index <= 7;
         when "0100111011010" => index <= 7;
         when "0100111011011" => index <= 6;
         when "0100111011100" => index <= 7;
         when "0100111011101" => index <= 6;
         when "0100111011110" => index <= 6;
         when "0100111011111" => index <= 6;
         when "0100111100000" => index <= 8;
         when "0100111100001" => index <= 7;
         when "0100111100010" => index <= 7;
         when "0100111100011" => index <= 6;
         when "0100111100100" => index <= 8;
         when "0100111100101" => index <= 7;
         when "0100111100110" => index <= 7;
         when "0100111100111" => index <= 6;
         when "0100111101000" => index <= 8;
         when "0100111101001" => index <= 7;
         when "0100111101010" => index <= 7;
         when "0100111101011" => index <= 6;
         when "0100111101100" => index <= 7;
         when "0100111101101" => index <= 6;
         when "0100111101110" => index <= 6;
         when "0100111101111" => index <= 6;
         when "0100111110000" => index <= 8;
         when "0100111110001" => index <= 7;
         when "0100111110010" => index <= 7;
         when "0100111110011" => index <= 6;
         when "0100111110100" => index <= 7;
         when "0100111110101" => index <= 6;
         when "0100111110110" => index <= 6;
         when "0100111110111" => index <= 6;
         when "0100111111000" => index <= 7;
         when "0100111111001" => index <= 6;
         when "0100111111010" => index <= 7;
         when "0100111111011" => index <= 6;
         when "0100111111100" => index <= 7;
         when "0100111111101" => index <= 6;
         when "0100111111110" => index <= 6;
         when "0100111111111" => index <= 6;
         when "0101000000000" => index <= 11;
         when "0101000000001" => index <= 8;
         when "0101000000010" => index <= 8;
         when "0101000000011" => index <= 6;
         when "0101000000100" => index <= 8;
         when "0101000000101" => index <= 6;
         when "0101000000110" => index <= 7;
         when "0101000000111" => index <= 6;
         when "0101000001000" => index <= 9;
         when "0101000001001" => index <= 7;
         when "0101000001010" => index <= 7;
         when "0101000001011" => index <= 6;
         when "0101000001100" => index <= 7;
         when "0101000001101" => index <= 6;
         when "0101000001110" => index <= 6;
         when "0101000001111" => index <= 5;
         when "0101000010000" => index <= 9;
         when "0101000010001" => index <= 7;
         when "0101000010010" => index <= 7;
         when "0101000010011" => index <= 6;
         when "0101000010100" => index <= 8;
         when "0101000010101" => index <= 6;
         when "0101000010110" => index <= 6;
         when "0101000010111" => index <= 6;
         when "0101000011000" => index <= 8;
         when "0101000011001" => index <= 6;
         when "0101000011010" => index <= 7;
         when "0101000011011" => index <= 6;
         when "0101000011100" => index <= 7;
         when "0101000011101" => index <= 6;
         when "0101000011110" => index <= 6;
         when "0101000011111" => index <= 5;
         when "0101000100000" => index <= 9;
         when "0101000100001" => index <= 7;
         when "0101000100010" => index <= 8;
         when "0101000100011" => index <= 6;
         when "0101000100100" => index <= 8;
         when "0101000100101" => index <= 6;
         when "0101000100110" => index <= 7;
         when "0101000100111" => index <= 6;
         when "0101000101000" => index <= 8;
         when "0101000101001" => index <= 7;
         when "0101000101010" => index <= 7;
         when "0101000101011" => index <= 6;
         when "0101000101100" => index <= 7;
         when "0101000101101" => index <= 6;
         when "0101000101110" => index <= 6;
         when "0101000101111" => index <= 5;
         when "0101000110000" => index <= 8;
         when "0101000110001" => index <= 7;
         when "0101000110010" => index <= 7;
         when "0101000110011" => index <= 6;
         when "0101000110100" => index <= 7;
         when "0101000110101" => index <= 6;
         when "0101000110110" => index <= 6;
         when "0101000110111" => index <= 6;
         when "0101000111000" => index <= 7;
         when "0101000111001" => index <= 6;
         when "0101000111010" => index <= 6;
         when "0101000111011" => index <= 6;
         when "0101000111100" => index <= 7;
         when "0101000111101" => index <= 6;
         when "0101000111110" => index <= 6;
         when "0101000111111" => index <= 5;
         when "0101001000000" => index <= 10;
         when "0101001000001" => index <= 8;
         when "0101001000010" => index <= 8;
         when "0101001000011" => index <= 6;
         when "0101001000100" => index <= 8;
         when "0101001000101" => index <= 7;
         when "0101001000110" => index <= 7;
         when "0101001000111" => index <= 6;
         when "0101001001000" => index <= 8;
         when "0101001001001" => index <= 7;
         when "0101001001010" => index <= 7;
         when "0101001001011" => index <= 6;
         when "0101001001100" => index <= 7;
         when "0101001001101" => index <= 6;
         when "0101001001110" => index <= 6;
         when "0101001001111" => index <= 6;
         when "0101001010000" => index <= 8;
         when "0101001010001" => index <= 7;
         when "0101001010010" => index <= 7;
         when "0101001010011" => index <= 6;
         when "0101001010100" => index <= 7;
         when "0101001010101" => index <= 6;
         when "0101001010110" => index <= 6;
         when "0101001010111" => index <= 6;
         when "0101001011000" => index <= 8;
         when "0101001011001" => index <= 6;
         when "0101001011010" => index <= 7;
         when "0101001011011" => index <= 6;
         when "0101001011100" => index <= 7;
         when "0101001011101" => index <= 6;
         when "0101001011110" => index <= 6;
         when "0101001011111" => index <= 6;
         when "0101001100000" => index <= 9;
         when "0101001100001" => index <= 7;
         when "0101001100010" => index <= 7;
         when "0101001100011" => index <= 6;
         when "0101001100100" => index <= 8;
         when "0101001100101" => index <= 6;
         when "0101001100110" => index <= 7;
         when "0101001100111" => index <= 6;
         when "0101001101000" => index <= 8;
         when "0101001101001" => index <= 7;
         when "0101001101010" => index <= 7;
         when "0101001101011" => index <= 6;
         when "0101001101100" => index <= 7;
         when "0101001101101" => index <= 6;
         when "0101001101110" => index <= 6;
         when "0101001101111" => index <= 6;
         when "0101001110000" => index <= 8;
         when "0101001110001" => index <= 7;
         when "0101001110010" => index <= 7;
         when "0101001110011" => index <= 6;
         when "0101001110100" => index <= 7;
         when "0101001110101" => index <= 6;
         when "0101001110110" => index <= 6;
         when "0101001110111" => index <= 6;
         when "0101001111000" => index <= 7;
         when "0101001111001" => index <= 6;
         when "0101001111010" => index <= 7;
         when "0101001111011" => index <= 6;
         when "0101001111100" => index <= 7;
         when "0101001111101" => index <= 6;
         when "0101001111110" => index <= 6;
         when "0101001111111" => index <= 6;
         when "0101010000000" => index <= 10;
         when "0101010000001" => index <= 8;
         when "0101010000010" => index <= 8;
         when "0101010000011" => index <= 7;
         when "0101010000100" => index <= 8;
         when "0101010000101" => index <= 7;
         when "0101010000110" => index <= 7;
         when "0101010000111" => index <= 6;
         when "0101010001000" => index <= 8;
         when "0101010001001" => index <= 7;
         when "0101010001010" => index <= 7;
         when "0101010001011" => index <= 6;
         when "0101010001100" => index <= 7;
         when "0101010001101" => index <= 6;
         when "0101010001110" => index <= 6;
         when "0101010001111" => index <= 6;
         when "0101010010000" => index <= 9;
         when "0101010010001" => index <= 7;
         when "0101010010010" => index <= 7;
         when "0101010010011" => index <= 6;
         when "0101010010100" => index <= 8;
         when "0101010010101" => index <= 6;
         when "0101010010110" => index <= 7;
         when "0101010010111" => index <= 6;
         when "0101010011000" => index <= 8;
         when "0101010011001" => index <= 7;
         when "0101010011010" => index <= 7;
         when "0101010011011" => index <= 6;
         when "0101010011100" => index <= 7;
         when "0101010011101" => index <= 6;
         when "0101010011110" => index <= 6;
         when "0101010011111" => index <= 6;
         when "0101010100000" => index <= 9;
         when "0101010100001" => index <= 7;
         when "0101010100010" => index <= 8;
         when "0101010100011" => index <= 6;
         when "0101010100100" => index <= 8;
         when "0101010100101" => index <= 7;
         when "0101010100110" => index <= 7;
         when "0101010100111" => index <= 6;
         when "0101010101000" => index <= 8;
         when "0101010101001" => index <= 7;
         when "0101010101010" => index <= 7;
         when "0101010101011" => index <= 6;
         when "0101010101100" => index <= 7;
         when "0101010101101" => index <= 6;
         when "0101010101110" => index <= 6;
         when "0101010101111" => index <= 6;
         when "0101010110000" => index <= 8;
         when "0101010110001" => index <= 7;
         when "0101010110010" => index <= 7;
         when "0101010110011" => index <= 6;
         when "0101010110100" => index <= 7;
         when "0101010110101" => index <= 6;
         when "0101010110110" => index <= 7;
         when "0101010110111" => index <= 6;
         when "0101010111000" => index <= 8;
         when "0101010111001" => index <= 7;
         when "0101010111010" => index <= 7;
         when "0101010111011" => index <= 6;
         when "0101010111100" => index <= 7;
         when "0101010111101" => index <= 6;
         when "0101010111110" => index <= 6;
         when "0101010111111" => index <= 6;
         when "0101011000000" => index <= 9;
         when "0101011000001" => index <= 8;
         when "0101011000010" => index <= 8;
         when "0101011000011" => index <= 7;
         when "0101011000100" => index <= 8;
         when "0101011000101" => index <= 7;
         when "0101011000110" => index <= 7;
         when "0101011000111" => index <= 6;
         when "0101011001000" => index <= 8;
         when "0101011001001" => index <= 7;
         when "0101011001010" => index <= 7;
         when "0101011001011" => index <= 6;
         when "0101011001100" => index <= 7;
         when "0101011001101" => index <= 6;
         when "0101011001110" => index <= 7;
         when "0101011001111" => index <= 6;
         when "0101011010000" => index <= 8;
         when "0101011010001" => index <= 7;
         when "0101011010010" => index <= 7;
         when "0101011010011" => index <= 6;
         when "0101011010100" => index <= 8;
         when "0101011010101" => index <= 7;
         when "0101011010110" => index <= 7;
         when "0101011010111" => index <= 6;
         when "0101011011000" => index <= 8;
         when "0101011011001" => index <= 7;
         when "0101011011010" => index <= 7;
         when "0101011011011" => index <= 6;
         when "0101011011100" => index <= 7;
         when "0101011011101" => index <= 6;
         when "0101011011110" => index <= 6;
         when "0101011011111" => index <= 6;
         when "0101011100000" => index <= 9;
         when "0101011100001" => index <= 7;
         when "0101011100010" => index <= 8;
         when "0101011100011" => index <= 7;
         when "0101011100100" => index <= 8;
         when "0101011100101" => index <= 7;
         when "0101011100110" => index <= 7;
         when "0101011100111" => index <= 6;
         when "0101011101000" => index <= 8;
         when "0101011101001" => index <= 7;
         when "0101011101010" => index <= 7;
         when "0101011101011" => index <= 6;
         when "0101011101100" => index <= 7;
         when "0101011101101" => index <= 6;
         when "0101011101110" => index <= 6;
         when "0101011101111" => index <= 6;
         when "0101011110000" => index <= 8;
         when "0101011110001" => index <= 7;
         when "0101011110010" => index <= 7;
         when "0101011110011" => index <= 6;
         when "0101011110100" => index <= 7;
         when "0101011110101" => index <= 6;
         when "0101011110110" => index <= 7;
         when "0101011110111" => index <= 6;
         when "0101011111000" => index <= 7;
         when "0101011111001" => index <= 7;
         when "0101011111010" => index <= 7;
         when "0101011111011" => index <= 6;
         when "0101011111100" => index <= 7;
         when "0101011111101" => index <= 6;
         when "0101011111110" => index <= 6;
         when "0101011111111" => index <= 6;
         when "0101100000000" => index <= 10;
         when "0101100000001" => index <= 8;
         when "0101100000010" => index <= 8;
         when "0101100000011" => index <= 7;
         when "0101100000100" => index <= 8;
         when "0101100000101" => index <= 7;
         when "0101100000110" => index <= 7;
         when "0101100000111" => index <= 6;
         when "0101100001000" => index <= 9;
         when "0101100001001" => index <= 7;
         when "0101100001010" => index <= 7;
         when "0101100001011" => index <= 6;
         when "0101100001100" => index <= 8;
         when "0101100001101" => index <= 6;
         when "0101100001110" => index <= 7;
         when "0101100001111" => index <= 6;
         when "0101100010000" => index <= 9;
         when "0101100010001" => index <= 7;
         when "0101100010010" => index <= 8;
         when "0101100010011" => index <= 6;
         when "0101100010100" => index <= 8;
         when "0101100010101" => index <= 7;
         when "0101100010110" => index <= 7;
         when "0101100010111" => index <= 6;
         when "0101100011000" => index <= 8;
         when "0101100011001" => index <= 7;
         when "0101100011010" => index <= 7;
         when "0101100011011" => index <= 6;
         when "0101100011100" => index <= 7;
         when "0101100011101" => index <= 6;
         when "0101100011110" => index <= 6;
         when "0101100011111" => index <= 6;
         when "0101100100000" => index <= 9;
         when "0101100100001" => index <= 8;
         when "0101100100010" => index <= 8;
         when "0101100100011" => index <= 7;
         when "0101100100100" => index <= 8;
         when "0101100100101" => index <= 7;
         when "0101100100110" => index <= 7;
         when "0101100100111" => index <= 6;
         when "0101100101000" => index <= 8;
         when "0101100101001" => index <= 7;
         when "0101100101010" => index <= 7;
         when "0101100101011" => index <= 6;
         when "0101100101100" => index <= 7;
         when "0101100101101" => index <= 6;
         when "0101100101110" => index <= 7;
         when "0101100101111" => index <= 6;
         when "0101100110000" => index <= 8;
         when "0101100110001" => index <= 7;
         when "0101100110010" => index <= 7;
         when "0101100110011" => index <= 6;
         when "0101100110100" => index <= 8;
         when "0101100110101" => index <= 7;
         when "0101100110110" => index <= 7;
         when "0101100110111" => index <= 6;
         when "0101100111000" => index <= 8;
         when "0101100111001" => index <= 7;
         when "0101100111010" => index <= 7;
         when "0101100111011" => index <= 6;
         when "0101100111100" => index <= 7;
         when "0101100111101" => index <= 6;
         when "0101100111110" => index <= 6;
         when "0101100111111" => index <= 6;
         when "0101101000000" => index <= 10;
         when "0101101000001" => index <= 8;
         when "0101101000010" => index <= 8;
         when "0101101000011" => index <= 7;
         when "0101101000100" => index <= 8;
         when "0101101000101" => index <= 7;
         when "0101101000110" => index <= 7;
         when "0101101000111" => index <= 6;
         when "0101101001000" => index <= 8;
         when "0101101001001" => index <= 7;
         when "0101101001010" => index <= 7;
         when "0101101001011" => index <= 6;
         when "0101101001100" => index <= 8;
         when "0101101001101" => index <= 7;
         when "0101101001110" => index <= 7;
         when "0101101001111" => index <= 6;
         when "0101101010000" => index <= 9;
         when "0101101010001" => index <= 7;
         when "0101101010010" => index <= 8;
         when "0101101010011" => index <= 7;
         when "0101101010100" => index <= 8;
         when "0101101010101" => index <= 7;
         when "0101101010110" => index <= 7;
         when "0101101010111" => index <= 6;
         when "0101101011000" => index <= 8;
         when "0101101011001" => index <= 7;
         when "0101101011010" => index <= 7;
         when "0101101011011" => index <= 6;
         when "0101101011100" => index <= 7;
         when "0101101011101" => index <= 6;
         when "0101101011110" => index <= 6;
         when "0101101011111" => index <= 6;
         when "0101101100000" => index <= 9;
         when "0101101100001" => index <= 8;
         when "0101101100010" => index <= 8;
         when "0101101100011" => index <= 7;
         when "0101101100100" => index <= 8;
         when "0101101100101" => index <= 7;
         when "0101101100110" => index <= 7;
         when "0101101100111" => index <= 6;
         when "0101101101000" => index <= 8;
         when "0101101101001" => index <= 7;
         when "0101101101010" => index <= 7;
         when "0101101101011" => index <= 6;
         when "0101101101100" => index <= 7;
         when "0101101101101" => index <= 6;
         when "0101101101110" => index <= 7;
         when "0101101101111" => index <= 6;
         when "0101101110000" => index <= 8;
         when "0101101110001" => index <= 7;
         when "0101101110010" => index <= 7;
         when "0101101110011" => index <= 6;
         when "0101101110100" => index <= 7;
         when "0101101110101" => index <= 7;
         when "0101101110110" => index <= 7;
         when "0101101110111" => index <= 6;
         when "0101101111000" => index <= 8;
         when "0101101111001" => index <= 7;
         when "0101101111010" => index <= 7;
         when "0101101111011" => index <= 6;
         when "0101101111100" => index <= 7;
         when "0101101111101" => index <= 6;
         when "0101101111110" => index <= 6;
         when "0101101111111" => index <= 6;
         when "0101110000000" => index <= 10;
         when "0101110000001" => index <= 8;
         when "0101110000010" => index <= 8;
         when "0101110000011" => index <= 7;
         when "0101110000100" => index <= 8;
         when "0101110000101" => index <= 7;
         when "0101110000110" => index <= 7;
         when "0101110000111" => index <= 6;
         when "0101110001000" => index <= 9;
         when "0101110001001" => index <= 7;
         when "0101110001010" => index <= 8;
         when "0101110001011" => index <= 7;
         when "0101110001100" => index <= 8;
         when "0101110001101" => index <= 7;
         when "0101110001110" => index <= 7;
         when "0101110001111" => index <= 6;
         when "0101110010000" => index <= 9;
         when "0101110010001" => index <= 8;
         when "0101110010010" => index <= 8;
         when "0101110010011" => index <= 7;
         when "0101110010100" => index <= 8;
         when "0101110010101" => index <= 7;
         when "0101110010110" => index <= 7;
         when "0101110010111" => index <= 6;
         when "0101110011000" => index <= 8;
         when "0101110011001" => index <= 7;
         when "0101110011010" => index <= 7;
         when "0101110011011" => index <= 6;
         when "0101110011100" => index <= 7;
         when "0101110011101" => index <= 6;
         when "0101110011110" => index <= 7;
         when "0101110011111" => index <= 6;
         when "0101110100000" => index <= 9;
         when "0101110100001" => index <= 8;
         when "0101110100010" => index <= 8;
         when "0101110100011" => index <= 7;
         when "0101110100100" => index <= 8;
         when "0101110100101" => index <= 7;
         when "0101110100110" => index <= 7;
         when "0101110100111" => index <= 6;
         when "0101110101000" => index <= 8;
         when "0101110101001" => index <= 7;
         when "0101110101010" => index <= 7;
         when "0101110101011" => index <= 6;
         when "0101110101100" => index <= 7;
         when "0101110101101" => index <= 7;
         when "0101110101110" => index <= 7;
         when "0101110101111" => index <= 6;
         when "0101110110000" => index <= 8;
         when "0101110110001" => index <= 7;
         when "0101110110010" => index <= 7;
         when "0101110110011" => index <= 7;
         when "0101110110100" => index <= 8;
         when "0101110110101" => index <= 7;
         when "0101110110110" => index <= 7;
         when "0101110110111" => index <= 6;
         when "0101110111000" => index <= 8;
         when "0101110111001" => index <= 7;
         when "0101110111010" => index <= 7;
         when "0101110111011" => index <= 6;
         when "0101110111100" => index <= 7;
         when "0101110111101" => index <= 6;
         when "0101110111110" => index <= 7;
         when "0101110111111" => index <= 6;
         when "0101111000000" => index <= 9;
         when "0101111000001" => index <= 8;
         when "0101111000010" => index <= 8;
         when "0101111000011" => index <= 7;
         when "0101111000100" => index <= 8;
         when "0101111000101" => index <= 7;
         when "0101111000110" => index <= 7;
         when "0101111000111" => index <= 6;
         when "0101111001000" => index <= 8;
         when "0101111001001" => index <= 7;
         when "0101111001010" => index <= 7;
         when "0101111001011" => index <= 7;
         when "0101111001100" => index <= 8;
         when "0101111001101" => index <= 7;
         when "0101111001110" => index <= 7;
         when "0101111001111" => index <= 6;
         when "0101111010000" => index <= 8;
         when "0101111010001" => index <= 7;
         when "0101111010010" => index <= 8;
         when "0101111010011" => index <= 7;
         when "0101111010100" => index <= 8;
         when "0101111010101" => index <= 7;
         when "0101111010110" => index <= 7;
         when "0101111010111" => index <= 6;
         when "0101111011000" => index <= 8;
         when "0101111011001" => index <= 7;
         when "0101111011010" => index <= 7;
         when "0101111011011" => index <= 6;
         when "0101111011100" => index <= 7;
         when "0101111011101" => index <= 7;
         when "0101111011110" => index <= 7;
         when "0101111011111" => index <= 6;
         when "0101111100000" => index <= 9;
         when "0101111100001" => index <= 8;
         when "0101111100010" => index <= 8;
         when "0101111100011" => index <= 7;
         when "0101111100100" => index <= 8;
         when "0101111100101" => index <= 7;
         when "0101111100110" => index <= 7;
         when "0101111100111" => index <= 6;
         when "0101111101000" => index <= 8;
         when "0101111101001" => index <= 7;
         when "0101111101010" => index <= 7;
         when "0101111101011" => index <= 7;
         when "0101111101100" => index <= 7;
         when "0101111101101" => index <= 7;
         when "0101111101110" => index <= 7;
         when "0101111101111" => index <= 6;
         when "0101111110000" => index <= 8;
         when "0101111110001" => index <= 7;
         when "0101111110010" => index <= 7;
         when "0101111110011" => index <= 7;
         when "0101111110100" => index <= 8;
         when "0101111110101" => index <= 7;
         when "0101111110110" => index <= 7;
         when "0101111110111" => index <= 6;
         when "0101111111000" => index <= 8;
         when "0101111111001" => index <= 7;
         when "0101111111010" => index <= 7;
         when "0101111111011" => index <= 6;
         when "0101111111100" => index <= 7;
         when "0101111111101" => index <= 6;
         when "0101111111110" => index <= 7;
         when "0101111111111" => index <= 6;
         when "0110000000000" => index <= 12;
         when "0110000000001" => index <= 8;
         when "0110000000010" => index <= 8;
         when "0110000000011" => index <= 6;
         when "0110000000100" => index <= 9;
         when "0110000000101" => index <= 7;
         when "0110000000110" => index <= 7;
         when "0110000000111" => index <= 6;
         when "0110000001000" => index <= 9;
         when "0110000001001" => index <= 7;
         when "0110000001010" => index <= 7;
         when "0110000001011" => index <= 6;
         when "0110000001100" => index <= 8;
         when "0110000001101" => index <= 6;
         when "0110000001110" => index <= 6;
         when "0110000001111" => index <= 6;
         when "0110000010000" => index <= 9;
         when "0110000010001" => index <= 7;
         when "0110000010010" => index <= 8;
         when "0110000010011" => index <= 6;
         when "0110000010100" => index <= 8;
         when "0110000010101" => index <= 6;
         when "0110000010110" => index <= 7;
         when "0110000010111" => index <= 6;
         when "0110000011000" => index <= 8;
         when "0110000011001" => index <= 7;
         when "0110000011010" => index <= 7;
         when "0110000011011" => index <= 6;
         when "0110000011100" => index <= 7;
         when "0110000011101" => index <= 6;
         when "0110000011110" => index <= 6;
         when "0110000011111" => index <= 5;
         when "0110000100000" => index <= 10;
         when "0110000100001" => index <= 8;
         when "0110000100010" => index <= 8;
         when "0110000100011" => index <= 6;
         when "0110000100100" => index <= 8;
         when "0110000100101" => index <= 7;
         when "0110000100110" => index <= 7;
         when "0110000100111" => index <= 6;
         when "0110000101000" => index <= 8;
         when "0110000101001" => index <= 7;
         when "0110000101010" => index <= 7;
         when "0110000101011" => index <= 6;
         when "0110000101100" => index <= 7;
         when "0110000101101" => index <= 6;
         when "0110000101110" => index <= 6;
         when "0110000101111" => index <= 6;
         when "0110000110000" => index <= 8;
         when "0110000110001" => index <= 7;
         when "0110000110010" => index <= 7;
         when "0110000110011" => index <= 6;
         when "0110000110100" => index <= 7;
         when "0110000110101" => index <= 6;
         when "0110000110110" => index <= 6;
         when "0110000110111" => index <= 6;
         when "0110000111000" => index <= 8;
         when "0110000111001" => index <= 6;
         when "0110000111010" => index <= 7;
         when "0110000111011" => index <= 6;
         when "0110000111100" => index <= 7;
         when "0110000111101" => index <= 6;
         when "0110000111110" => index <= 6;
         when "0110000111111" => index <= 6;
         when "0110001000000" => index <= 10;
         when "0110001000001" => index <= 8;
         when "0110001000010" => index <= 8;
         when "0110001000011" => index <= 7;
         when "0110001000100" => index <= 8;
         when "0110001000101" => index <= 7;
         when "0110001000110" => index <= 7;
         when "0110001000111" => index <= 6;
         when "0110001001000" => index <= 8;
         when "0110001001001" => index <= 7;
         when "0110001001010" => index <= 7;
         when "0110001001011" => index <= 6;
         when "0110001001100" => index <= 7;
         when "0110001001101" => index <= 6;
         when "0110001001110" => index <= 6;
         when "0110001001111" => index <= 6;
         when "0110001010000" => index <= 9;
         when "0110001010001" => index <= 7;
         when "0110001010010" => index <= 7;
         when "0110001010011" => index <= 6;
         when "0110001010100" => index <= 8;
         when "0110001010101" => index <= 6;
         when "0110001010110" => index <= 7;
         when "0110001010111" => index <= 6;
         when "0110001011000" => index <= 8;
         when "0110001011001" => index <= 7;
         when "0110001011010" => index <= 7;
         when "0110001011011" => index <= 6;
         when "0110001011100" => index <= 7;
         when "0110001011101" => index <= 6;
         when "0110001011110" => index <= 6;
         when "0110001011111" => index <= 6;
         when "0110001100000" => index <= 9;
         when "0110001100001" => index <= 7;
         when "0110001100010" => index <= 8;
         when "0110001100011" => index <= 6;
         when "0110001100100" => index <= 8;
         when "0110001100101" => index <= 7;
         when "0110001100110" => index <= 7;
         when "0110001100111" => index <= 6;
         when "0110001101000" => index <= 8;
         when "0110001101001" => index <= 7;
         when "0110001101010" => index <= 7;
         when "0110001101011" => index <= 6;
         when "0110001101100" => index <= 7;
         when "0110001101101" => index <= 6;
         when "0110001101110" => index <= 6;
         when "0110001101111" => index <= 6;
         when "0110001110000" => index <= 8;
         when "0110001110001" => index <= 7;
         when "0110001110010" => index <= 7;
         when "0110001110011" => index <= 6;
         when "0110001110100" => index <= 7;
         when "0110001110101" => index <= 6;
         when "0110001110110" => index <= 7;
         when "0110001110111" => index <= 6;
         when "0110001111000" => index <= 8;
         when "0110001111001" => index <= 7;
         when "0110001111010" => index <= 7;
         when "0110001111011" => index <= 6;
         when "0110001111100" => index <= 7;
         when "0110001111101" => index <= 6;
         when "0110001111110" => index <= 6;
         when "0110001111111" => index <= 6;
         when "0110010000000" => index <= 10;
         when "0110010000001" => index <= 8;
         when "0110010000010" => index <= 8;
         when "0110010000011" => index <= 7;
         when "0110010000100" => index <= 8;
         when "0110010000101" => index <= 7;
         when "0110010000110" => index <= 7;
         when "0110010000111" => index <= 6;
         when "0110010001000" => index <= 9;
         when "0110010001001" => index <= 7;
         when "0110010001010" => index <= 7;
         when "0110010001011" => index <= 6;
         when "0110010001100" => index <= 8;
         when "0110010001101" => index <= 6;
         when "0110010001110" => index <= 7;
         when "0110010001111" => index <= 6;
         when "0110010010000" => index <= 9;
         when "0110010010001" => index <= 7;
         when "0110010010010" => index <= 8;
         when "0110010010011" => index <= 6;
         when "0110010010100" => index <= 8;
         when "0110010010101" => index <= 7;
         when "0110010010110" => index <= 7;
         when "0110010010111" => index <= 6;
         when "0110010011000" => index <= 8;
         when "0110010011001" => index <= 7;
         when "0110010011010" => index <= 7;
         when "0110010011011" => index <= 6;
         when "0110010011100" => index <= 7;
         when "0110010011101" => index <= 6;
         when "0110010011110" => index <= 6;
         when "0110010011111" => index <= 6;
         when "0110010100000" => index <= 9;
         when "0110010100001" => index <= 8;
         when "0110010100010" => index <= 8;
         when "0110010100011" => index <= 7;
         when "0110010100100" => index <= 8;
         when "0110010100101" => index <= 7;
         when "0110010100110" => index <= 7;
         when "0110010100111" => index <= 6;
         when "0110010101000" => index <= 8;
         when "0110010101001" => index <= 7;
         when "0110010101010" => index <= 7;
         when "0110010101011" => index <= 6;
         when "0110010101100" => index <= 7;
         when "0110010101101" => index <= 6;
         when "0110010101110" => index <= 7;
         when "0110010101111" => index <= 6;
         when "0110010110000" => index <= 8;
         when "0110010110001" => index <= 7;
         when "0110010110010" => index <= 7;
         when "0110010110011" => index <= 6;
         when "0110010110100" => index <= 8;
         when "0110010110101" => index <= 7;
         when "0110010110110" => index <= 7;
         when "0110010110111" => index <= 6;
         when "0110010111000" => index <= 8;
         when "0110010111001" => index <= 7;
         when "0110010111010" => index <= 7;
         when "0110010111011" => index <= 6;
         when "0110010111100" => index <= 7;
         when "0110010111101" => index <= 6;
         when "0110010111110" => index <= 6;
         when "0110010111111" => index <= 6;
         when "0110011000000" => index <= 10;
         when "0110011000001" => index <= 8;
         when "0110011000010" => index <= 8;
         when "0110011000011" => index <= 7;
         when "0110011000100" => index <= 8;
         when "0110011000101" => index <= 7;
         when "0110011000110" => index <= 7;
         when "0110011000111" => index <= 6;
         when "0110011001000" => index <= 8;
         when "0110011001001" => index <= 7;
         when "0110011001010" => index <= 7;
         when "0110011001011" => index <= 6;
         when "0110011001100" => index <= 8;
         when "0110011001101" => index <= 7;
         when "0110011001110" => index <= 7;
         when "0110011001111" => index <= 6;
         when "0110011010000" => index <= 9;
         when "0110011010001" => index <= 7;
         when "0110011010010" => index <= 8;
         when "0110011010011" => index <= 7;
         when "0110011010100" => index <= 8;
         when "0110011010101" => index <= 7;
         when "0110011010110" => index <= 7;
         when "0110011010111" => index <= 6;
         when "0110011011000" => index <= 8;
         when "0110011011001" => index <= 7;
         when "0110011011010" => index <= 7;
         when "0110011011011" => index <= 6;
         when "0110011011100" => index <= 7;
         when "0110011011101" => index <= 6;
         when "0110011011110" => index <= 6;
         when "0110011011111" => index <= 6;
         when "0110011100000" => index <= 9;
         when "0110011100001" => index <= 8;
         when "0110011100010" => index <= 8;
         when "0110011100011" => index <= 7;
         when "0110011100100" => index <= 8;
         when "0110011100101" => index <= 7;
         when "0110011100110" => index <= 7;
         when "0110011100111" => index <= 6;
         when "0110011101000" => index <= 8;
         when "0110011101001" => index <= 7;
         when "0110011101010" => index <= 7;
         when "0110011101011" => index <= 6;
         when "0110011101100" => index <= 7;
         when "0110011101101" => index <= 6;
         when "0110011101110" => index <= 7;
         when "0110011101111" => index <= 6;
         when "0110011110000" => index <= 8;
         when "0110011110001" => index <= 7;
         when "0110011110010" => index <= 7;
         when "0110011110011" => index <= 6;
         when "0110011110100" => index <= 7;
         when "0110011110101" => index <= 7;
         when "0110011110110" => index <= 7;
         when "0110011110111" => index <= 6;
         when "0110011111000" => index <= 8;
         when "0110011111001" => index <= 7;
         when "0110011111010" => index <= 7;
         when "0110011111011" => index <= 6;
         when "0110011111100" => index <= 7;
         when "0110011111101" => index <= 6;
         when "0110011111110" => index <= 6;
         when "0110011111111" => index <= 6;
         when "0110100000000" => index <= 11;
         when "0110100000001" => index <= 8;
         when "0110100000010" => index <= 8;
         when "0110100000011" => index <= 7;
         when "0110100000100" => index <= 9;
         when "0110100000101" => index <= 7;
         when "0110100000110" => index <= 7;
         when "0110100000111" => index <= 6;
         when "0110100001000" => index <= 9;
         when "0110100001001" => index <= 7;
         when "0110100001010" => index <= 8;
         when "0110100001011" => index <= 6;
         when "0110100001100" => index <= 8;
         when "0110100001101" => index <= 7;
         when "0110100001110" => index <= 7;
         when "0110100001111" => index <= 6;
         when "0110100010000" => index <= 9;
         when "0110100010001" => index <= 8;
         when "0110100010010" => index <= 8;
         when "0110100010011" => index <= 7;
         when "0110100010100" => index <= 8;
         when "0110100010101" => index <= 7;
         when "0110100010110" => index <= 7;
         when "0110100010111" => index <= 6;
         when "0110100011000" => index <= 8;
         when "0110100011001" => index <= 7;
         when "0110100011010" => index <= 7;
         when "0110100011011" => index <= 6;
         when "0110100011100" => index <= 7;
         when "0110100011101" => index <= 6;
         when "0110100011110" => index <= 7;
         when "0110100011111" => index <= 6;
         when "0110100100000" => index <= 10;
         when "0110100100001" => index <= 8;
         when "0110100100010" => index <= 8;
         when "0110100100011" => index <= 7;
         when "0110100100100" => index <= 8;
         when "0110100100101" => index <= 7;
         when "0110100100110" => index <= 7;
         when "0110100100111" => index <= 6;
         when "0110100101000" => index <= 8;
         when "0110100101001" => index <= 7;
         when "0110100101010" => index <= 7;
         when "0110100101011" => index <= 6;
         when "0110100101100" => index <= 8;
         when "0110100101101" => index <= 7;
         when "0110100101110" => index <= 7;
         when "0110100101111" => index <= 6;
         when "0110100110000" => index <= 9;
         when "0110100110001" => index <= 7;
         when "0110100110010" => index <= 8;
         when "0110100110011" => index <= 7;
         when "0110100110100" => index <= 8;
         when "0110100110101" => index <= 7;
         when "0110100110110" => index <= 7;
         when "0110100110111" => index <= 6;
         when "0110100111000" => index <= 8;
         when "0110100111001" => index <= 7;
         when "0110100111010" => index <= 7;
         when "0110100111011" => index <= 6;
         when "0110100111100" => index <= 7;
         when "0110100111101" => index <= 6;
         when "0110100111110" => index <= 6;
         when "0110100111111" => index <= 6;
         when "0110101000000" => index <= 10;
         when "0110101000001" => index <= 8;
         when "0110101000010" => index <= 8;
         when "0110101000011" => index <= 7;
         when "0110101000100" => index <= 8;
         when "0110101000101" => index <= 7;
         when "0110101000110" => index <= 7;
         when "0110101000111" => index <= 6;
         when "0110101001000" => index <= 9;
         when "0110101001001" => index <= 7;
         when "0110101001010" => index <= 8;
         when "0110101001011" => index <= 7;
         when "0110101001100" => index <= 8;
         when "0110101001101" => index <= 7;
         when "0110101001110" => index <= 7;
         when "0110101001111" => index <= 6;
         when "0110101010000" => index <= 9;
         when "0110101010001" => index <= 8;
         when "0110101010010" => index <= 8;
         when "0110101010011" => index <= 7;
         when "0110101010100" => index <= 8;
         when "0110101010101" => index <= 7;
         when "0110101010110" => index <= 7;
         when "0110101010111" => index <= 6;
         when "0110101011000" => index <= 8;
         when "0110101011001" => index <= 7;
         when "0110101011010" => index <= 7;
         when "0110101011011" => index <= 6;
         when "0110101011100" => index <= 7;
         when "0110101011101" => index <= 6;
         when "0110101011110" => index <= 7;
         when "0110101011111" => index <= 6;
         when "0110101100000" => index <= 9;
         when "0110101100001" => index <= 8;
         when "0110101100010" => index <= 8;
         when "0110101100011" => index <= 7;
         when "0110101100100" => index <= 8;
         when "0110101100101" => index <= 7;
         when "0110101100110" => index <= 7;
         when "0110101100111" => index <= 6;
         when "0110101101000" => index <= 8;
         when "0110101101001" => index <= 7;
         when "0110101101010" => index <= 7;
         when "0110101101011" => index <= 6;
         when "0110101101100" => index <= 7;
         when "0110101101101" => index <= 7;
         when "0110101101110" => index <= 7;
         when "0110101101111" => index <= 6;
         when "0110101110000" => index <= 8;
         when "0110101110001" => index <= 7;
         when "0110101110010" => index <= 7;
         when "0110101110011" => index <= 7;
         when "0110101110100" => index <= 8;
         when "0110101110101" => index <= 7;
         when "0110101110110" => index <= 7;
         when "0110101110111" => index <= 6;
         when "0110101111000" => index <= 8;
         when "0110101111001" => index <= 7;
         when "0110101111010" => index <= 7;
         when "0110101111011" => index <= 6;
         when "0110101111100" => index <= 7;
         when "0110101111101" => index <= 6;
         when "0110101111110" => index <= 7;
         when "0110101111111" => index <= 6;
         when "0110110000000" => index <= 10;
         when "0110110000001" => index <= 8;
         when "0110110000010" => index <= 8;
         when "0110110000011" => index <= 7;
         when "0110110000100" => index <= 9;
         when "0110110000101" => index <= 7;
         when "0110110000110" => index <= 8;
         when "0110110000111" => index <= 7;
         when "0110110001000" => index <= 9;
         when "0110110001001" => index <= 8;
         when "0110110001010" => index <= 8;
         when "0110110001011" => index <= 7;
         when "0110110001100" => index <= 8;
         when "0110110001101" => index <= 7;
         when "0110110001110" => index <= 7;
         when "0110110001111" => index <= 6;
         when "0110110010000" => index <= 9;
         when "0110110010001" => index <= 8;
         when "0110110010010" => index <= 8;
         when "0110110010011" => index <= 7;
         when "0110110010100" => index <= 8;
         when "0110110010101" => index <= 7;
         when "0110110010110" => index <= 7;
         when "0110110010111" => index <= 6;
         when "0110110011000" => index <= 8;
         when "0110110011001" => index <= 7;
         when "0110110011010" => index <= 7;
         when "0110110011011" => index <= 6;
         when "0110110011100" => index <= 7;
         when "0110110011101" => index <= 7;
         when "0110110011110" => index <= 7;
         when "0110110011111" => index <= 6;
         when "0110110100000" => index <= 9;
         when "0110110100001" => index <= 8;
         when "0110110100010" => index <= 8;
         when "0110110100011" => index <= 7;
         when "0110110100100" => index <= 8;
         when "0110110100101" => index <= 7;
         when "0110110100110" => index <= 7;
         when "0110110100111" => index <= 6;
         when "0110110101000" => index <= 8;
         when "0110110101001" => index <= 7;
         when "0110110101010" => index <= 7;
         when "0110110101011" => index <= 7;
         when "0110110101100" => index <= 8;
         when "0110110101101" => index <= 7;
         when "0110110101110" => index <= 7;
         when "0110110101111" => index <= 6;
         when "0110110110000" => index <= 8;
         when "0110110110001" => index <= 7;
         when "0110110110010" => index <= 8;
         when "0110110110011" => index <= 7;
         when "0110110110100" => index <= 8;
         when "0110110110101" => index <= 7;
         when "0110110110110" => index <= 7;
         when "0110110110111" => index <= 6;
         when "0110110111000" => index <= 8;
         when "0110110111001" => index <= 7;
         when "0110110111010" => index <= 7;
         when "0110110111011" => index <= 6;
         when "0110110111100" => index <= 7;
         when "0110110111101" => index <= 7;
         when "0110110111110" => index <= 7;
         when "0110110111111" => index <= 6;
         when "0110111000000" => index <= 9;
         when "0110111000001" => index <= 8;
         when "0110111000010" => index <= 8;
         when "0110111000011" => index <= 7;
         when "0110111000100" => index <= 8;
         when "0110111000101" => index <= 7;
         when "0110111000110" => index <= 7;
         when "0110111000111" => index <= 7;
         when "0110111001000" => index <= 8;
         when "0110111001001" => index <= 7;
         when "0110111001010" => index <= 8;
         when "0110111001011" => index <= 7;
         when "0110111001100" => index <= 8;
         when "0110111001101" => index <= 7;
         when "0110111001110" => index <= 7;
         when "0110111001111" => index <= 6;
         when "0110111010000" => index <= 9;
         when "0110111010001" => index <= 8;
         when "0110111010010" => index <= 8;
         when "0110111010011" => index <= 7;
         when "0110111010100" => index <= 8;
         when "0110111010101" => index <= 7;
         when "0110111010110" => index <= 7;
         when "0110111010111" => index <= 6;
         when "0110111011000" => index <= 8;
         when "0110111011001" => index <= 7;
         when "0110111011010" => index <= 7;
         when "0110111011011" => index <= 7;
         when "0110111011100" => index <= 7;
         when "0110111011101" => index <= 7;
         when "0110111011110" => index <= 7;
         when "0110111011111" => index <= 6;
         when "0110111100000" => index <= 9;
         when "0110111100001" => index <= 8;
         when "0110111100010" => index <= 8;
         when "0110111100011" => index <= 7;
         when "0110111100100" => index <= 8;
         when "0110111100101" => index <= 7;
         when "0110111100110" => index <= 7;
         when "0110111100111" => index <= 7;
         when "0110111101000" => index <= 8;
         when "0110111101001" => index <= 7;
         when "0110111101010" => index <= 7;
         when "0110111101011" => index <= 7;
         when "0110111101100" => index <= 8;
         when "0110111101101" => index <= 7;
         when "0110111101110" => index <= 7;
         when "0110111101111" => index <= 6;
         when "0110111110000" => index <= 8;
         when "0110111110001" => index <= 7;
         when "0110111110010" => index <= 8;
         when "0110111110011" => index <= 7;
         when "0110111110100" => index <= 8;
         when "0110111110101" => index <= 7;
         when "0110111110110" => index <= 7;
         when "0110111110111" => index <= 6;
         when "0110111111000" => index <= 8;
         when "0110111111001" => index <= 7;
         when "0110111111010" => index <= 7;
         when "0110111111011" => index <= 6;
         when "0110111111100" => index <= 7;
         when "0110111111101" => index <= 7;
         when "0110111111110" => index <= 7;
         when "0110111111111" => index <= 6;
         when "0111000000000" => index <= 11;
         when "0111000000001" => index <= 8;
         when "0111000000010" => index <= 9;
         when "0111000000011" => index <= 7;
         when "0111000000100" => index <= 9;
         when "0111000000101" => index <= 7;
         when "0111000000110" => index <= 8;
         when "0111000000111" => index <= 6;
         when "0111000001000" => index <= 9;
         when "0111000001001" => index <= 8;
         when "0111000001010" => index <= 8;
         when "0111000001011" => index <= 7;
         when "0111000001100" => index <= 8;
         when "0111000001101" => index <= 7;
         when "0111000001110" => index <= 7;
         when "0111000001111" => index <= 6;
         when "0111000010000" => index <= 10;
         when "0111000010001" => index <= 8;
         when "0111000010010" => index <= 8;
         when "0111000010011" => index <= 7;
         when "0111000010100" => index <= 8;
         when "0111000010101" => index <= 7;
         when "0111000010110" => index <= 7;
         when "0111000010111" => index <= 6;
         when "0111000011000" => index <= 8;
         when "0111000011001" => index <= 7;
         when "0111000011010" => index <= 7;
         when "0111000011011" => index <= 6;
         when "0111000011100" => index <= 8;
         when "0111000011101" => index <= 7;
         when "0111000011110" => index <= 7;
         when "0111000011111" => index <= 6;
         when "0111000100000" => index <= 10;
         when "0111000100001" => index <= 8;
         when "0111000100010" => index <= 8;
         when "0111000100011" => index <= 7;
         when "0111000100100" => index <= 8;
         when "0111000100101" => index <= 7;
         when "0111000100110" => index <= 7;
         when "0111000100111" => index <= 6;
         when "0111000101000" => index <= 9;
         when "0111000101001" => index <= 7;
         when "0111000101010" => index <= 8;
         when "0111000101011" => index <= 7;
         when "0111000101100" => index <= 8;
         when "0111000101101" => index <= 7;
         when "0111000101110" => index <= 7;
         when "0111000101111" => index <= 6;
         when "0111000110000" => index <= 9;
         when "0111000110001" => index <= 8;
         when "0111000110010" => index <= 8;
         when "0111000110011" => index <= 7;
         when "0111000110100" => index <= 8;
         when "0111000110101" => index <= 7;
         when "0111000110110" => index <= 7;
         when "0111000110111" => index <= 6;
         when "0111000111000" => index <= 8;
         when "0111000111001" => index <= 7;
         when "0111000111010" => index <= 7;
         when "0111000111011" => index <= 6;
         when "0111000111100" => index <= 7;
         when "0111000111101" => index <= 6;
         when "0111000111110" => index <= 7;
         when "0111000111111" => index <= 6;
         when "0111001000000" => index <= 10;
         when "0111001000001" => index <= 8;
         when "0111001000010" => index <= 8;
         when "0111001000011" => index <= 7;
         when "0111001000100" => index <= 9;
         when "0111001000101" => index <= 7;
         when "0111001000110" => index <= 8;
         when "0111001000111" => index <= 7;
         when "0111001001000" => index <= 9;
         when "0111001001001" => index <= 8;
         when "0111001001010" => index <= 8;
         when "0111001001011" => index <= 7;
         when "0111001001100" => index <= 8;
         when "0111001001101" => index <= 7;
         when "0111001001110" => index <= 7;
         when "0111001001111" => index <= 6;
         when "0111001010000" => index <= 9;
         when "0111001010001" => index <= 8;
         when "0111001010010" => index <= 8;
         when "0111001010011" => index <= 7;
         when "0111001010100" => index <= 8;
         when "0111001010101" => index <= 7;
         when "0111001010110" => index <= 7;
         when "0111001010111" => index <= 6;
         when "0111001011000" => index <= 8;
         when "0111001011001" => index <= 7;
         when "0111001011010" => index <= 7;
         when "0111001011011" => index <= 6;
         when "0111001011100" => index <= 7;
         when "0111001011101" => index <= 7;
         when "0111001011110" => index <= 7;
         when "0111001011111" => index <= 6;
         when "0111001100000" => index <= 9;
         when "0111001100001" => index <= 8;
         when "0111001100010" => index <= 8;
         when "0111001100011" => index <= 7;
         when "0111001100100" => index <= 8;
         when "0111001100101" => index <= 7;
         when "0111001100110" => index <= 7;
         when "0111001100111" => index <= 6;
         when "0111001101000" => index <= 8;
         when "0111001101001" => index <= 7;
         when "0111001101010" => index <= 7;
         when "0111001101011" => index <= 7;
         when "0111001101100" => index <= 8;
         when "0111001101101" => index <= 7;
         when "0111001101110" => index <= 7;
         when "0111001101111" => index <= 6;
         when "0111001110000" => index <= 8;
         when "0111001110001" => index <= 7;
         when "0111001110010" => index <= 8;
         when "0111001110011" => index <= 7;
         when "0111001110100" => index <= 8;
         when "0111001110101" => index <= 7;
         when "0111001110110" => index <= 7;
         when "0111001110111" => index <= 6;
         when "0111001111000" => index <= 8;
         when "0111001111001" => index <= 7;
         when "0111001111010" => index <= 7;
         when "0111001111011" => index <= 6;
         when "0111001111100" => index <= 7;
         when "0111001111101" => index <= 7;
         when "0111001111110" => index <= 7;
         when "0111001111111" => index <= 6;
         when "0111010000000" => index <= 10;
         when "0111010000001" => index <= 8;
         when "0111010000010" => index <= 9;
         when "0111010000011" => index <= 7;
         when "0111010000100" => index <= 9;
         when "0111010000101" => index <= 8;
         when "0111010000110" => index <= 8;
         when "0111010000111" => index <= 7;
         when "0111010001000" => index <= 9;
         when "0111010001001" => index <= 8;
         when "0111010001010" => index <= 8;
         when "0111010001011" => index <= 7;
         when "0111010001100" => index <= 8;
         when "0111010001101" => index <= 7;
         when "0111010001110" => index <= 7;
         when "0111010001111" => index <= 6;
         when "0111010010000" => index <= 9;
         when "0111010010001" => index <= 8;
         when "0111010010010" => index <= 8;
         when "0111010010011" => index <= 7;
         when "0111010010100" => index <= 8;
         when "0111010010101" => index <= 7;
         when "0111010010110" => index <= 7;
         when "0111010010111" => index <= 6;
         when "0111010011000" => index <= 8;
         when "0111010011001" => index <= 7;
         when "0111010011010" => index <= 7;
         when "0111010011011" => index <= 7;
         when "0111010011100" => index <= 8;
         when "0111010011101" => index <= 7;
         when "0111010011110" => index <= 7;
         when "0111010011111" => index <= 6;
         when "0111010100000" => index <= 9;
         when "0111010100001" => index <= 8;
         when "0111010100010" => index <= 8;
         when "0111010100011" => index <= 7;
         when "0111010100100" => index <= 8;
         when "0111010100101" => index <= 7;
         when "0111010100110" => index <= 7;
         when "0111010100111" => index <= 7;
         when "0111010101000" => index <= 8;
         when "0111010101001" => index <= 7;
         when "0111010101010" => index <= 8;
         when "0111010101011" => index <= 7;
         when "0111010101100" => index <= 8;
         when "0111010101101" => index <= 7;
         when "0111010101110" => index <= 7;
         when "0111010101111" => index <= 6;
         when "0111010110000" => index <= 9;
         when "0111010110001" => index <= 8;
         when "0111010110010" => index <= 8;
         when "0111010110011" => index <= 7;
         when "0111010110100" => index <= 8;
         when "0111010110101" => index <= 7;
         when "0111010110110" => index <= 7;
         when "0111010110111" => index <= 6;
         when "0111010111000" => index <= 8;
         when "0111010111001" => index <= 7;
         when "0111010111010" => index <= 7;
         when "0111010111011" => index <= 7;
         when "0111010111100" => index <= 7;
         when "0111010111101" => index <= 7;
         when "0111010111110" => index <= 7;
         when "0111010111111" => index <= 6;
         when "0111011000000" => index <= 10;
         when "0111011000001" => index <= 8;
         when "0111011000010" => index <= 8;
         when "0111011000011" => index <= 7;
         when "0111011000100" => index <= 8;
         when "0111011000101" => index <= 7;
         when "0111011000110" => index <= 8;
         when "0111011000111" => index <= 7;
         when "0111011001000" => index <= 9;
         when "0111011001001" => index <= 8;
         when "0111011001010" => index <= 8;
         when "0111011001011" => index <= 7;
         when "0111011001100" => index <= 8;
         when "0111011001101" => index <= 7;
         when "0111011001110" => index <= 7;
         when "0111011001111" => index <= 6;
         when "0111011010000" => index <= 9;
         when "0111011010001" => index <= 8;
         when "0111011010010" => index <= 8;
         when "0111011010011" => index <= 7;
         when "0111011010100" => index <= 8;
         when "0111011010101" => index <= 7;
         when "0111011010110" => index <= 7;
         when "0111011010111" => index <= 7;
         when "0111011011000" => index <= 8;
         when "0111011011001" => index <= 7;
         when "0111011011010" => index <= 7;
         when "0111011011011" => index <= 7;
         when "0111011011100" => index <= 8;
         when "0111011011101" => index <= 7;
         when "0111011011110" => index <= 7;
         when "0111011011111" => index <= 6;
         when "0111011100000" => index <= 9;
         when "0111011100001" => index <= 8;
         when "0111011100010" => index <= 8;
         when "0111011100011" => index <= 7;
         when "0111011100100" => index <= 8;
         when "0111011100101" => index <= 7;
         when "0111011100110" => index <= 7;
         when "0111011100111" => index <= 7;
         when "0111011101000" => index <= 8;
         when "0111011101001" => index <= 7;
         when "0111011101010" => index <= 8;
         when "0111011101011" => index <= 7;
         when "0111011101100" => index <= 8;
         when "0111011101101" => index <= 7;
         when "0111011101110" => index <= 7;
         when "0111011101111" => index <= 6;
         when "0111011110000" => index <= 8;
         when "0111011110001" => index <= 8;
         when "0111011110010" => index <= 8;
         when "0111011110011" => index <= 7;
         when "0111011110100" => index <= 8;
         when "0111011110101" => index <= 7;
         when "0111011110110" => index <= 7;
         when "0111011110111" => index <= 6;
         when "0111011111000" => index <= 8;
         when "0111011111001" => index <= 7;
         when "0111011111010" => index <= 7;
         when "0111011111011" => index <= 7;
         when "0111011111100" => index <= 7;
         when "0111011111101" => index <= 7;
         when "0111011111110" => index <= 7;
         when "0111011111111" => index <= 6;
         when "0111100000000" => index <= 10;
         when "0111100000001" => index <= 9;
         when "0111100000010" => index <= 9;
         when "0111100000011" => index <= 8;
         when "0111100000100" => index <= 9;
         when "0111100000101" => index <= 8;
         when "0111100000110" => index <= 8;
         when "0111100000111" => index <= 7;
         when "0111100001000" => index <= 9;
         when "0111100001001" => index <= 8;
         when "0111100001010" => index <= 8;
         when "0111100001011" => index <= 7;
         when "0111100001100" => index <= 8;
         when "0111100001101" => index <= 7;
         when "0111100001110" => index <= 7;
         when "0111100001111" => index <= 6;
         when "0111100010000" => index <= 9;
         when "0111100010001" => index <= 8;
         when "0111100010010" => index <= 8;
         when "0111100010011" => index <= 7;
         when "0111100010100" => index <= 8;
         when "0111100010101" => index <= 7;
         when "0111100010110" => index <= 7;
         when "0111100010111" => index <= 7;
         when "0111100011000" => index <= 8;
         when "0111100011001" => index <= 7;
         when "0111100011010" => index <= 8;
         when "0111100011011" => index <= 7;
         when "0111100011100" => index <= 8;
         when "0111100011101" => index <= 7;
         when "0111100011110" => index <= 7;
         when "0111100011111" => index <= 6;
         when "0111100100000" => index <= 10;
         when "0111100100001" => index <= 8;
         when "0111100100010" => index <= 8;
         when "0111100100011" => index <= 7;
         when "0111100100100" => index <= 8;
         when "0111100100101" => index <= 7;
         when "0111100100110" => index <= 8;
         when "0111100100111" => index <= 7;
         when "0111100101000" => index <= 9;
         when "0111100101001" => index <= 8;
         when "0111100101010" => index <= 8;
         when "0111100101011" => index <= 7;
         when "0111100101100" => index <= 8;
         when "0111100101101" => index <= 7;
         when "0111100101110" => index <= 7;
         when "0111100101111" => index <= 6;
         when "0111100110000" => index <= 9;
         when "0111100110001" => index <= 8;
         when "0111100110010" => index <= 8;
         when "0111100110011" => index <= 7;
         when "0111100110100" => index <= 8;
         when "0111100110101" => index <= 7;
         when "0111100110110" => index <= 7;
         when "0111100110111" => index <= 7;
         when "0111100111000" => index <= 8;
         when "0111100111001" => index <= 7;
         when "0111100111010" => index <= 7;
         when "0111100111011" => index <= 7;
         when "0111100111100" => index <= 8;
         when "0111100111101" => index <= 7;
         when "0111100111110" => index <= 7;
         when "0111100111111" => index <= 6;
         when "0111101000000" => index <= 10;
         when "0111101000001" => index <= 8;
         when "0111101000010" => index <= 8;
         when "0111101000011" => index <= 7;
         when "0111101000100" => index <= 9;
         when "0111101000101" => index <= 8;
         when "0111101000110" => index <= 8;
         when "0111101000111" => index <= 7;
         when "0111101001000" => index <= 9;
         when "0111101001001" => index <= 8;
         when "0111101001010" => index <= 8;
         when "0111101001011" => index <= 7;
         when "0111101001100" => index <= 8;
         when "0111101001101" => index <= 7;
         when "0111101001110" => index <= 7;
         when "0111101001111" => index <= 7;
         when "0111101010000" => index <= 9;
         when "0111101010001" => index <= 8;
         when "0111101010010" => index <= 8;
         when "0111101010011" => index <= 7;
         when "0111101010100" => index <= 8;
         when "0111101010101" => index <= 7;
         when "0111101010110" => index <= 7;
         when "0111101010111" => index <= 7;
         when "0111101011000" => index <= 8;
         when "0111101011001" => index <= 7;
         when "0111101011010" => index <= 8;
         when "0111101011011" => index <= 7;
         when "0111101011100" => index <= 8;
         when "0111101011101" => index <= 7;
         when "0111101011110" => index <= 7;
         when "0111101011111" => index <= 6;
         when "0111101100000" => index <= 9;
         when "0111101100001" => index <= 8;
         when "0111101100010" => index <= 8;
         when "0111101100011" => index <= 7;
         when "0111101100100" => index <= 8;
         when "0111101100101" => index <= 7;
         when "0111101100110" => index <= 8;
         when "0111101100111" => index <= 7;
         when "0111101101000" => index <= 8;
         when "0111101101001" => index <= 8;
         when "0111101101010" => index <= 8;
         when "0111101101011" => index <= 7;
         when "0111101101100" => index <= 8;
         when "0111101101101" => index <= 7;
         when "0111101101110" => index <= 7;
         when "0111101101111" => index <= 6;
         when "0111101110000" => index <= 9;
         when "0111101110001" => index <= 8;
         when "0111101110010" => index <= 8;
         when "0111101110011" => index <= 7;
         when "0111101110100" => index <= 8;
         when "0111101110101" => index <= 7;
         when "0111101110110" => index <= 7;
         when "0111101110111" => index <= 7;
         when "0111101111000" => index <= 8;
         when "0111101111001" => index <= 7;
         when "0111101111010" => index <= 7;
         when "0111101111011" => index <= 7;
         when "0111101111100" => index <= 7;
         when "0111101111101" => index <= 7;
         when "0111101111110" => index <= 7;
         when "0111101111111" => index <= 6;
         when "0111110000000" => index <= 10;
         when "0111110000001" => index <= 8;
         when "0111110000010" => index <= 9;
         when "0111110000011" => index <= 8;
         when "0111110000100" => index <= 9;
         when "0111110000101" => index <= 8;
         when "0111110000110" => index <= 8;
         when "0111110000111" => index <= 7;
         when "0111110001000" => index <= 9;
         when "0111110001001" => index <= 8;
         when "0111110001010" => index <= 8;
         when "0111110001011" => index <= 7;
         when "0111110001100" => index <= 8;
         when "0111110001101" => index <= 7;
         when "0111110001110" => index <= 7;
         when "0111110001111" => index <= 7;
         when "0111110010000" => index <= 9;
         when "0111110010001" => index <= 8;
         when "0111110010010" => index <= 8;
         when "0111110010011" => index <= 7;
         when "0111110010100" => index <= 8;
         when "0111110010101" => index <= 7;
         when "0111110010110" => index <= 8;
         when "0111110010111" => index <= 7;
         when "0111110011000" => index <= 8;
         when "0111110011001" => index <= 8;
         when "0111110011010" => index <= 8;
         when "0111110011011" => index <= 7;
         when "0111110011100" => index <= 8;
         when "0111110011101" => index <= 7;
         when "0111110011110" => index <= 7;
         when "0111110011111" => index <= 6;
         when "0111110100000" => index <= 9;
         when "0111110100001" => index <= 8;
         when "0111110100010" => index <= 8;
         when "0111110100011" => index <= 7;
         when "0111110100100" => index <= 8;
         when "0111110100101" => index <= 8;
         when "0111110100110" => index <= 8;
         when "0111110100111" => index <= 7;
         when "0111110101000" => index <= 9;
         when "0111110101001" => index <= 8;
         when "0111110101010" => index <= 8;
         when "0111110101011" => index <= 7;
         when "0111110101100" => index <= 8;
         when "0111110101101" => index <= 7;
         when "0111110101110" => index <= 7;
         when "0111110101111" => index <= 7;
         when "0111110110000" => index <= 9;
         when "0111110110001" => index <= 8;
         when "0111110110010" => index <= 8;
         when "0111110110011" => index <= 7;
         when "0111110110100" => index <= 8;
         when "0111110110101" => index <= 7;
         when "0111110110110" => index <= 7;
         when "0111110110111" => index <= 7;
         when "0111110111000" => index <= 8;
         when "0111110111001" => index <= 7;
         when "0111110111010" => index <= 7;
         when "0111110111011" => index <= 7;
         when "0111110111100" => index <= 8;
         when "0111110111101" => index <= 7;
         when "0111110111110" => index <= 7;
         when "0111110111111" => index <= 6;
         when "0111111000000" => index <= 10;
         when "0111111000001" => index <= 8;
         when "0111111000010" => index <= 8;
         when "0111111000011" => index <= 8;
         when "0111111000100" => index <= 9;
         when "0111111000101" => index <= 8;
         when "0111111000110" => index <= 8;
         when "0111111000111" => index <= 7;
         when "0111111001000" => index <= 9;
         when "0111111001001" => index <= 8;
         when "0111111001010" => index <= 8;
         when "0111111001011" => index <= 7;
         when "0111111001100" => index <= 8;
         when "0111111001101" => index <= 7;
         when "0111111001110" => index <= 7;
         when "0111111001111" => index <= 7;
         when "0111111010000" => index <= 9;
         when "0111111010001" => index <= 8;
         when "0111111010010" => index <= 8;
         when "0111111010011" => index <= 7;
         when "0111111010100" => index <= 8;
         when "0111111010101" => index <= 7;
         when "0111111010110" => index <= 7;
         when "0111111010111" => index <= 7;
         when "0111111011000" => index <= 8;
         when "0111111011001" => index <= 7;
         when "0111111011010" => index <= 8;
         when "0111111011011" => index <= 7;
         when "0111111011100" => index <= 8;
         when "0111111011101" => index <= 7;
         when "0111111011110" => index <= 7;
         when "0111111011111" => index <= 7;
         when "0111111100000" => index <= 9;
         when "0111111100001" => index <= 8;
         when "0111111100010" => index <= 8;
         when "0111111100011" => index <= 7;
         when "0111111100100" => index <= 8;
         when "0111111100101" => index <= 7;
         when "0111111100110" => index <= 8;
         when "0111111100111" => index <= 7;
         when "0111111101000" => index <= 8;
         when "0111111101001" => index <= 8;
         when "0111111101010" => index <= 8;
         when "0111111101011" => index <= 7;
         when "0111111101100" => index <= 8;
         when "0111111101101" => index <= 7;
         when "0111111101110" => index <= 7;
         when "0111111101111" => index <= 7;
         when "0111111110000" => index <= 8;
         when "0111111110001" => index <= 8;
         when "0111111110010" => index <= 8;
         when "0111111110011" => index <= 7;
         when "0111111110100" => index <= 8;
         when "0111111110101" => index <= 7;
         when "0111111110110" => index <= 7;
         when "0111111110111" => index <= 7;
         when "0111111111000" => index <= 8;
         when "0111111111001" => index <= 7;
         when "0111111111010" => index <= 7;
         when "0111111111011" => index <= 7;
         when "0111111111100" => index <= 8;
         when "0111111111101" => index <= 7;
         when "0111111111110" => index <= 7;
         when "0111111111111" => index <= 6;
         when "1000000000000" => index <= 13;
         when "1000000000001" => index <= 7;
         when "1000000000010" => index <= 8;
         when "1000000000011" => index <= 5;
         when "1000000000100" => index <= 8;
         when "1000000000101" => index <= 6;
         when "1000000000110" => index <= 6;
         when "1000000000111" => index <= 5;
         when "1000000001000" => index <= 8;
         when "1000000001001" => index <= 6;
         when "1000000001010" => index <= 6;
         when "1000000001011" => index <= 5;
         when "1000000001100" => index <= 7;
         when "1000000001101" => index <= 5;
         when "1000000001110" => index <= 6;
         when "1000000001111" => index <= 5;
         when "1000000010000" => index <= 9;
         when "1000000010001" => index <= 6;
         when "1000000010010" => index <= 7;
         when "1000000010011" => index <= 5;
         when "1000000010100" => index <= 7;
         when "1000000010101" => index <= 6;
         when "1000000010110" => index <= 6;
         when "1000000010111" => index <= 5;
         when "1000000011000" => index <= 7;
         when "1000000011001" => index <= 6;
         when "1000000011010" => index <= 6;
         when "1000000011011" => index <= 5;
         when "1000000011100" => index <= 6;
         when "1000000011101" => index <= 5;
         when "1000000011110" => index <= 5;
         when "1000000011111" => index <= 5;
         when "1000000100000" => index <= 10;
         when "1000000100001" => index <= 7;
         when "1000000100010" => index <= 7;
         when "1000000100011" => index <= 6;
         when "1000000100100" => index <= 7;
         when "1000000100101" => index <= 6;
         when "1000000100110" => index <= 6;
         when "1000000100111" => index <= 5;
         when "1000000101000" => index <= 8;
         when "1000000101001" => index <= 6;
         when "1000000101010" => index <= 6;
         when "1000000101011" => index <= 5;
         when "1000000101100" => index <= 6;
         when "1000000101101" => index <= 5;
         when "1000000101110" => index <= 6;
         when "1000000101111" => index <= 5;
         when "1000000110000" => index <= 8;
         when "1000000110001" => index <= 6;
         when "1000000110010" => index <= 6;
         when "1000000110011" => index <= 5;
         when "1000000110100" => index <= 7;
         when "1000000110101" => index <= 6;
         when "1000000110110" => index <= 6;
         when "1000000110111" => index <= 5;
         when "1000000111000" => index <= 7;
         when "1000000111001" => index <= 6;
         when "1000000111010" => index <= 6;
         when "1000000111011" => index <= 5;
         when "1000000111100" => index <= 6;
         when "1000000111101" => index <= 5;
         when "1000000111110" => index <= 6;
         when "1000000111111" => index <= 5;
         when "1000001000000" => index <= 10;
         when "1000001000001" => index <= 7;
         when "1000001000010" => index <= 7;
         when "1000001000011" => index <= 6;
         when "1000001000100" => index <= 8;
         when "1000001000101" => index <= 6;
         when "1000001000110" => index <= 6;
         when "1000001000111" => index <= 5;
         when "1000001001000" => index <= 8;
         when "1000001001001" => index <= 6;
         when "1000001001010" => index <= 6;
         when "1000001001011" => index <= 5;
         when "1000001001100" => index <= 7;
         when "1000001001101" => index <= 6;
         when "1000001001110" => index <= 6;
         when "1000001001111" => index <= 5;
         when "1000001010000" => index <= 8;
         when "1000001010001" => index <= 6;
         when "1000001010010" => index <= 7;
         when "1000001010011" => index <= 6;
         when "1000001010100" => index <= 7;
         when "1000001010101" => index <= 6;
         when "1000001010110" => index <= 6;
         when "1000001010111" => index <= 5;
         when "1000001011000" => index <= 7;
         when "1000001011001" => index <= 6;
         when "1000001011010" => index <= 6;
         when "1000001011011" => index <= 5;
         when "1000001011100" => index <= 6;
         when "1000001011101" => index <= 6;
         when "1000001011110" => index <= 6;
         when "1000001011111" => index <= 5;
         when "1000001100000" => index <= 9;
         when "1000001100001" => index <= 7;
         when "1000001100010" => index <= 7;
         when "1000001100011" => index <= 6;
         when "1000001100100" => index <= 7;
         when "1000001100101" => index <= 6;
         when "1000001100110" => index <= 6;
         when "1000001100111" => index <= 5;
         when "1000001101000" => index <= 8;
         when "1000001101001" => index <= 6;
         when "1000001101010" => index <= 6;
         when "1000001101011" => index <= 6;
         when "1000001101100" => index <= 7;
         when "1000001101101" => index <= 6;
         when "1000001101110" => index <= 6;
         when "1000001101111" => index <= 5;
         when "1000001110000" => index <= 8;
         when "1000001110001" => index <= 6;
         when "1000001110010" => index <= 7;
         when "1000001110011" => index <= 6;
         when "1000001110100" => index <= 7;
         when "1000001110101" => index <= 6;
         when "1000001110110" => index <= 6;
         when "1000001110111" => index <= 5;
         when "1000001111000" => index <= 7;
         when "1000001111001" => index <= 6;
         when "1000001111010" => index <= 6;
         when "1000001111011" => index <= 5;
         when "1000001111100" => index <= 6;
         when "1000001111101" => index <= 6;
         when "1000001111110" => index <= 6;
         when "1000001111111" => index <= 5;
         when "1000010000000" => index <= 10;
         when "1000010000001" => index <= 7;
         when "1000010000010" => index <= 8;
         when "1000010000011" => index <= 6;
         when "1000010000100" => index <= 8;
         when "1000010000101" => index <= 6;
         when "1000010000110" => index <= 6;
         when "1000010000111" => index <= 5;
         when "1000010001000" => index <= 8;
         when "1000010001001" => index <= 6;
         when "1000010001010" => index <= 7;
         when "1000010001011" => index <= 6;
         when "1000010001100" => index <= 7;
         when "1000010001101" => index <= 6;
         when "1000010001110" => index <= 6;
         when "1000010001111" => index <= 5;
         when "1000010010000" => index <= 9;
         when "1000010010001" => index <= 7;
         when "1000010010010" => index <= 7;
         when "1000010010011" => index <= 6;
         when "1000010010100" => index <= 7;
         when "1000010010101" => index <= 6;
         when "1000010010110" => index <= 6;
         when "1000010010111" => index <= 5;
         when "1000010011000" => index <= 8;
         when "1000010011001" => index <= 6;
         when "1000010011010" => index <= 6;
         when "1000010011011" => index <= 6;
         when "1000010011100" => index <= 7;
         when "1000010011101" => index <= 6;
         when "1000010011110" => index <= 6;
         when "1000010011111" => index <= 5;
         when "1000010100000" => index <= 9;
         when "1000010100001" => index <= 7;
         when "1000010100010" => index <= 7;
         when "1000010100011" => index <= 6;
         when "1000010100100" => index <= 8;
         when "1000010100101" => index <= 6;
         when "1000010100110" => index <= 6;
         when "1000010100111" => index <= 6;
         when "1000010101000" => index <= 8;
         when "1000010101001" => index <= 6;
         when "1000010101010" => index <= 7;
         when "1000010101011" => index <= 6;
         when "1000010101100" => index <= 7;
         when "1000010101101" => index <= 6;
         when "1000010101110" => index <= 6;
         when "1000010101111" => index <= 5;
         when "1000010110000" => index <= 8;
         when "1000010110001" => index <= 7;
         when "1000010110010" => index <= 7;
         when "1000010110011" => index <= 6;
         when "1000010110100" => index <= 7;
         when "1000010110101" => index <= 6;
         when "1000010110110" => index <= 6;
         when "1000010110111" => index <= 5;
         when "1000010111000" => index <= 7;
         when "1000010111001" => index <= 6;
         when "1000010111010" => index <= 6;
         when "1000010111011" => index <= 6;
         when "1000010111100" => index <= 6;
         when "1000010111101" => index <= 6;
         when "1000010111110" => index <= 6;
         when "1000010111111" => index <= 5;
         when "1000011000000" => index <= 9;
         when "1000011000001" => index <= 7;
         when "1000011000010" => index <= 8;
         when "1000011000011" => index <= 6;
         when "1000011000100" => index <= 8;
         when "1000011000101" => index <= 6;
         when "1000011000110" => index <= 7;
         when "1000011000111" => index <= 6;
         when "1000011001000" => index <= 8;
         when "1000011001001" => index <= 7;
         when "1000011001010" => index <= 7;
         when "1000011001011" => index <= 6;
         when "1000011001100" => index <= 7;
         when "1000011001101" => index <= 6;
         when "1000011001110" => index <= 6;
         when "1000011001111" => index <= 5;
         when "1000011010000" => index <= 8;
         when "1000011010001" => index <= 7;
         when "1000011010010" => index <= 7;
         when "1000011010011" => index <= 6;
         when "1000011010100" => index <= 7;
         when "1000011010101" => index <= 6;
         when "1000011010110" => index <= 6;
         when "1000011010111" => index <= 6;
         when "1000011011000" => index <= 7;
         when "1000011011001" => index <= 6;
         when "1000011011010" => index <= 6;
         when "1000011011011" => index <= 6;
         when "1000011011100" => index <= 7;
         when "1000011011101" => index <= 6;
         when "1000011011110" => index <= 6;
         when "1000011011111" => index <= 5;
         when "1000011100000" => index <= 8;
         when "1000011100001" => index <= 7;
         when "1000011100010" => index <= 7;
         when "1000011100011" => index <= 6;
         when "1000011100100" => index <= 7;
         when "1000011100101" => index <= 6;
         when "1000011100110" => index <= 6;
         when "1000011100111" => index <= 6;
         when "1000011101000" => index <= 8;
         when "1000011101001" => index <= 6;
         when "1000011101010" => index <= 7;
         when "1000011101011" => index <= 6;
         when "1000011101100" => index <= 7;
         when "1000011101101" => index <= 6;
         when "1000011101110" => index <= 6;
         when "1000011101111" => index <= 6;
         when "1000011110000" => index <= 8;
         when "1000011110001" => index <= 7;
         when "1000011110010" => index <= 7;
         when "1000011110011" => index <= 6;
         when "1000011110100" => index <= 7;
         when "1000011110101" => index <= 6;
         when "1000011110110" => index <= 6;
         when "1000011110111" => index <= 6;
         when "1000011111000" => index <= 7;
         when "1000011111001" => index <= 6;
         when "1000011111010" => index <= 6;
         when "1000011111011" => index <= 6;
         when "1000011111100" => index <= 7;
         when "1000011111101" => index <= 6;
         when "1000011111110" => index <= 6;
         when "1000011111111" => index <= 5;
         when "1000100000000" => index <= 11;
         when "1000100000001" => index <= 8;
         when "1000100000010" => index <= 8;
         when "1000100000011" => index <= 6;
         when "1000100000100" => index <= 8;
         when "1000100000101" => index <= 6;
         when "1000100000110" => index <= 7;
         when "1000100000111" => index <= 6;
         when "1000100001000" => index <= 9;
         when "1000100001001" => index <= 7;
         when "1000100001010" => index <= 7;
         when "1000100001011" => index <= 6;
         when "1000100001100" => index <= 7;
         when "1000100001101" => index <= 6;
         when "1000100001110" => index <= 6;
         when "1000100001111" => index <= 5;
         when "1000100010000" => index <= 9;
         when "1000100010001" => index <= 7;
         when "1000100010010" => index <= 7;
         when "1000100010011" => index <= 6;
         when "1000100010100" => index <= 8;
         when "1000100010101" => index <= 6;
         when "1000100010110" => index <= 6;
         when "1000100010111" => index <= 6;
         when "1000100011000" => index <= 8;
         when "1000100011001" => index <= 6;
         when "1000100011010" => index <= 7;
         when "1000100011011" => index <= 6;
         when "1000100011100" => index <= 7;
         when "1000100011101" => index <= 6;
         when "1000100011110" => index <= 6;
         when "1000100011111" => index <= 5;
         when "1000100100000" => index <= 9;
         when "1000100100001" => index <= 7;
         when "1000100100010" => index <= 8;
         when "1000100100011" => index <= 6;
         when "1000100100100" => index <= 8;
         when "1000100100101" => index <= 6;
         when "1000100100110" => index <= 7;
         when "1000100100111" => index <= 6;
         when "1000100101000" => index <= 8;
         when "1000100101001" => index <= 7;
         when "1000100101010" => index <= 7;
         when "1000100101011" => index <= 6;
         when "1000100101100" => index <= 7;
         when "1000100101101" => index <= 6;
         when "1000100101110" => index <= 6;
         when "1000100101111" => index <= 5;
         when "1000100110000" => index <= 8;
         when "1000100110001" => index <= 7;
         when "1000100110010" => index <= 7;
         when "1000100110011" => index <= 6;
         when "1000100110100" => index <= 7;
         when "1000100110101" => index <= 6;
         when "1000100110110" => index <= 6;
         when "1000100110111" => index <= 6;
         when "1000100111000" => index <= 7;
         when "1000100111001" => index <= 6;
         when "1000100111010" => index <= 6;
         when "1000100111011" => index <= 6;
         when "1000100111100" => index <= 7;
         when "1000100111101" => index <= 6;
         when "1000100111110" => index <= 6;
         when "1000100111111" => index <= 5;
         when "1000101000000" => index <= 10;
         when "1000101000001" => index <= 8;
         when "1000101000010" => index <= 8;
         when "1000101000011" => index <= 6;
         when "1000101000100" => index <= 8;
         when "1000101000101" => index <= 7;
         when "1000101000110" => index <= 7;
         when "1000101000111" => index <= 6;
         when "1000101001000" => index <= 8;
         when "1000101001001" => index <= 7;
         when "1000101001010" => index <= 7;
         when "1000101001011" => index <= 6;
         when "1000101001100" => index <= 7;
         when "1000101001101" => index <= 6;
         when "1000101001110" => index <= 6;
         when "1000101001111" => index <= 6;
         when "1000101010000" => index <= 8;
         when "1000101010001" => index <= 7;
         when "1000101010010" => index <= 7;
         when "1000101010011" => index <= 6;
         when "1000101010100" => index <= 7;
         when "1000101010101" => index <= 6;
         when "1000101010110" => index <= 6;
         when "1000101010111" => index <= 6;
         when "1000101011000" => index <= 8;
         when "1000101011001" => index <= 6;
         when "1000101011010" => index <= 7;
         when "1000101011011" => index <= 6;
         when "1000101011100" => index <= 7;
         when "1000101011101" => index <= 6;
         when "1000101011110" => index <= 6;
         when "1000101011111" => index <= 6;
         when "1000101100000" => index <= 9;
         when "1000101100001" => index <= 7;
         when "1000101100010" => index <= 7;
         when "1000101100011" => index <= 6;
         when "1000101100100" => index <= 8;
         when "1000101100101" => index <= 6;
         when "1000101100110" => index <= 7;
         when "1000101100111" => index <= 6;
         when "1000101101000" => index <= 8;
         when "1000101101001" => index <= 7;
         when "1000101101010" => index <= 7;
         when "1000101101011" => index <= 6;
         when "1000101101100" => index <= 7;
         when "1000101101101" => index <= 6;
         when "1000101101110" => index <= 6;
         when "1000101101111" => index <= 6;
         when "1000101110000" => index <= 8;
         when "1000101110001" => index <= 7;
         when "1000101110010" => index <= 7;
         when "1000101110011" => index <= 6;
         when "1000101110100" => index <= 7;
         when "1000101110101" => index <= 6;
         when "1000101110110" => index <= 6;
         when "1000101110111" => index <= 6;
         when "1000101111000" => index <= 7;
         when "1000101111001" => index <= 6;
         when "1000101111010" => index <= 7;
         when "1000101111011" => index <= 6;
         when "1000101111100" => index <= 7;
         when "1000101111101" => index <= 6;
         when "1000101111110" => index <= 6;
         when "1000101111111" => index <= 6;
         when "1000110000000" => index <= 10;
         when "1000110000001" => index <= 8;
         when "1000110000010" => index <= 8;
         when "1000110000011" => index <= 7;
         when "1000110000100" => index <= 8;
         when "1000110000101" => index <= 7;
         when "1000110000110" => index <= 7;
         when "1000110000111" => index <= 6;
         when "1000110001000" => index <= 8;
         when "1000110001001" => index <= 7;
         when "1000110001010" => index <= 7;
         when "1000110001011" => index <= 6;
         when "1000110001100" => index <= 7;
         when "1000110001101" => index <= 6;
         when "1000110001110" => index <= 6;
         when "1000110001111" => index <= 6;
         when "1000110010000" => index <= 9;
         when "1000110010001" => index <= 7;
         when "1000110010010" => index <= 7;
         when "1000110010011" => index <= 6;
         when "1000110010100" => index <= 8;
         when "1000110010101" => index <= 6;
         when "1000110010110" => index <= 7;
         when "1000110010111" => index <= 6;
         when "1000110011000" => index <= 8;
         when "1000110011001" => index <= 7;
         when "1000110011010" => index <= 7;
         when "1000110011011" => index <= 6;
         when "1000110011100" => index <= 7;
         when "1000110011101" => index <= 6;
         when "1000110011110" => index <= 6;
         when "1000110011111" => index <= 6;
         when "1000110100000" => index <= 9;
         when "1000110100001" => index <= 7;
         when "1000110100010" => index <= 8;
         when "1000110100011" => index <= 6;
         when "1000110100100" => index <= 8;
         when "1000110100101" => index <= 7;
         when "1000110100110" => index <= 7;
         when "1000110100111" => index <= 6;
         when "1000110101000" => index <= 8;
         when "1000110101001" => index <= 7;
         when "1000110101010" => index <= 7;
         when "1000110101011" => index <= 6;
         when "1000110101100" => index <= 7;
         when "1000110101101" => index <= 6;
         when "1000110101110" => index <= 6;
         when "1000110101111" => index <= 6;
         when "1000110110000" => index <= 8;
         when "1000110110001" => index <= 7;
         when "1000110110010" => index <= 7;
         when "1000110110011" => index <= 6;
         when "1000110110100" => index <= 7;
         when "1000110110101" => index <= 6;
         when "1000110110110" => index <= 7;
         when "1000110110111" => index <= 6;
         when "1000110111000" => index <= 8;
         when "1000110111001" => index <= 7;
         when "1000110111010" => index <= 7;
         when "1000110111011" => index <= 6;
         when "1000110111100" => index <= 7;
         when "1000110111101" => index <= 6;
         when "1000110111110" => index <= 6;
         when "1000110111111" => index <= 6;
         when "1000111000000" => index <= 9;
         when "1000111000001" => index <= 8;
         when "1000111000010" => index <= 8;
         when "1000111000011" => index <= 7;
         when "1000111000100" => index <= 8;
         when "1000111000101" => index <= 7;
         when "1000111000110" => index <= 7;
         when "1000111000111" => index <= 6;
         when "1000111001000" => index <= 8;
         when "1000111001001" => index <= 7;
         when "1000111001010" => index <= 7;
         when "1000111001011" => index <= 6;
         when "1000111001100" => index <= 7;
         when "1000111001101" => index <= 6;
         when "1000111001110" => index <= 7;
         when "1000111001111" => index <= 6;
         when "1000111010000" => index <= 8;
         when "1000111010001" => index <= 7;
         when "1000111010010" => index <= 7;
         when "1000111010011" => index <= 6;
         when "1000111010100" => index <= 8;
         when "1000111010101" => index <= 7;
         when "1000111010110" => index <= 7;
         when "1000111010111" => index <= 6;
         when "1000111011000" => index <= 8;
         when "1000111011001" => index <= 7;
         when "1000111011010" => index <= 7;
         when "1000111011011" => index <= 6;
         when "1000111011100" => index <= 7;
         when "1000111011101" => index <= 6;
         when "1000111011110" => index <= 6;
         when "1000111011111" => index <= 6;
         when "1000111100000" => index <= 9;
         when "1000111100001" => index <= 7;
         when "1000111100010" => index <= 8;
         when "1000111100011" => index <= 7;
         when "1000111100100" => index <= 8;
         when "1000111100101" => index <= 7;
         when "1000111100110" => index <= 7;
         when "1000111100111" => index <= 6;
         when "1000111101000" => index <= 8;
         when "1000111101001" => index <= 7;
         when "1000111101010" => index <= 7;
         when "1000111101011" => index <= 6;
         when "1000111101100" => index <= 7;
         when "1000111101101" => index <= 6;
         when "1000111101110" => index <= 6;
         when "1000111101111" => index <= 6;
         when "1000111110000" => index <= 8;
         when "1000111110001" => index <= 7;
         when "1000111110010" => index <= 7;
         when "1000111110011" => index <= 6;
         when "1000111110100" => index <= 7;
         when "1000111110101" => index <= 6;
         when "1000111110110" => index <= 7;
         when "1000111110111" => index <= 6;
         when "1000111111000" => index <= 7;
         when "1000111111001" => index <= 7;
         when "1000111111010" => index <= 7;
         when "1000111111011" => index <= 6;
         when "1000111111100" => index <= 7;
         when "1000111111101" => index <= 6;
         when "1000111111110" => index <= 6;
         when "1000111111111" => index <= 6;
         when "1001000000000" => index <= 12;
         when "1001000000001" => index <= 8;
         when "1001000000010" => index <= 8;
         when "1001000000011" => index <= 6;
         when "1001000000100" => index <= 9;
         when "1001000000101" => index <= 7;
         when "1001000000110" => index <= 7;
         when "1001000000111" => index <= 6;
         when "1001000001000" => index <= 9;
         when "1001000001001" => index <= 7;
         when "1001000001010" => index <= 7;
         when "1001000001011" => index <= 6;
         when "1001000001100" => index <= 8;
         when "1001000001101" => index <= 6;
         when "1001000001110" => index <= 6;
         when "1001000001111" => index <= 6;
         when "1001000010000" => index <= 9;
         when "1001000010001" => index <= 7;
         when "1001000010010" => index <= 8;
         when "1001000010011" => index <= 6;
         when "1001000010100" => index <= 8;
         when "1001000010101" => index <= 6;
         when "1001000010110" => index <= 7;
         when "1001000010111" => index <= 6;
         when "1001000011000" => index <= 8;
         when "1001000011001" => index <= 7;
         when "1001000011010" => index <= 7;
         when "1001000011011" => index <= 6;
         when "1001000011100" => index <= 7;
         when "1001000011101" => index <= 6;
         when "1001000011110" => index <= 6;
         when "1001000011111" => index <= 5;
         when "1001000100000" => index <= 10;
         when "1001000100001" => index <= 8;
         when "1001000100010" => index <= 8;
         when "1001000100011" => index <= 6;
         when "1001000100100" => index <= 8;
         when "1001000100101" => index <= 7;
         when "1001000100110" => index <= 7;
         when "1001000100111" => index <= 6;
         when "1001000101000" => index <= 8;
         when "1001000101001" => index <= 7;
         when "1001000101010" => index <= 7;
         when "1001000101011" => index <= 6;
         when "1001000101100" => index <= 7;
         when "1001000101101" => index <= 6;
         when "1001000101110" => index <= 6;
         when "1001000101111" => index <= 6;
         when "1001000110000" => index <= 8;
         when "1001000110001" => index <= 7;
         when "1001000110010" => index <= 7;
         when "1001000110011" => index <= 6;
         when "1001000110100" => index <= 7;
         when "1001000110101" => index <= 6;
         when "1001000110110" => index <= 6;
         when "1001000110111" => index <= 6;
         when "1001000111000" => index <= 8;
         when "1001000111001" => index <= 6;
         when "1001000111010" => index <= 7;
         when "1001000111011" => index <= 6;
         when "1001000111100" => index <= 7;
         when "1001000111101" => index <= 6;
         when "1001000111110" => index <= 6;
         when "1001000111111" => index <= 6;
         when "1001001000000" => index <= 10;
         when "1001001000001" => index <= 8;
         when "1001001000010" => index <= 8;
         when "1001001000011" => index <= 7;
         when "1001001000100" => index <= 8;
         when "1001001000101" => index <= 7;
         when "1001001000110" => index <= 7;
         when "1001001000111" => index <= 6;
         when "1001001001000" => index <= 8;
         when "1001001001001" => index <= 7;
         when "1001001001010" => index <= 7;
         when "1001001001011" => index <= 6;
         when "1001001001100" => index <= 7;
         when "1001001001101" => index <= 6;
         when "1001001001110" => index <= 6;
         when "1001001001111" => index <= 6;
         when "1001001010000" => index <= 9;
         when "1001001010001" => index <= 7;
         when "1001001010010" => index <= 7;
         when "1001001010011" => index <= 6;
         when "1001001010100" => index <= 8;
         when "1001001010101" => index <= 6;
         when "1001001010110" => index <= 7;
         when "1001001010111" => index <= 6;
         when "1001001011000" => index <= 8;
         when "1001001011001" => index <= 7;
         when "1001001011010" => index <= 7;
         when "1001001011011" => index <= 6;
         when "1001001011100" => index <= 7;
         when "1001001011101" => index <= 6;
         when "1001001011110" => index <= 6;
         when "1001001011111" => index <= 6;
         when "1001001100000" => index <= 9;
         when "1001001100001" => index <= 7;
         when "1001001100010" => index <= 8;
         when "1001001100011" => index <= 6;
         when "1001001100100" => index <= 8;
         when "1001001100101" => index <= 7;
         when "1001001100110" => index <= 7;
         when "1001001100111" => index <= 6;
         when "1001001101000" => index <= 8;
         when "1001001101001" => index <= 7;
         when "1001001101010" => index <= 7;
         when "1001001101011" => index <= 6;
         when "1001001101100" => index <= 7;
         when "1001001101101" => index <= 6;
         when "1001001101110" => index <= 6;
         when "1001001101111" => index <= 6;
         when "1001001110000" => index <= 8;
         when "1001001110001" => index <= 7;
         when "1001001110010" => index <= 7;
         when "1001001110011" => index <= 6;
         when "1001001110100" => index <= 7;
         when "1001001110101" => index <= 6;
         when "1001001110110" => index <= 7;
         when "1001001110111" => index <= 6;
         when "1001001111000" => index <= 8;
         when "1001001111001" => index <= 7;
         when "1001001111010" => index <= 7;
         when "1001001111011" => index <= 6;
         when "1001001111100" => index <= 7;
         when "1001001111101" => index <= 6;
         when "1001001111110" => index <= 6;
         when "1001001111111" => index <= 6;
         when "1001010000000" => index <= 10;
         when "1001010000001" => index <= 8;
         when "1001010000010" => index <= 8;
         when "1001010000011" => index <= 7;
         when "1001010000100" => index <= 8;
         when "1001010000101" => index <= 7;
         when "1001010000110" => index <= 7;
         when "1001010000111" => index <= 6;
         when "1001010001000" => index <= 9;
         when "1001010001001" => index <= 7;
         when "1001010001010" => index <= 7;
         when "1001010001011" => index <= 6;
         when "1001010001100" => index <= 8;
         when "1001010001101" => index <= 6;
         when "1001010001110" => index <= 7;
         when "1001010001111" => index <= 6;
         when "1001010010000" => index <= 9;
         when "1001010010001" => index <= 7;
         when "1001010010010" => index <= 8;
         when "1001010010011" => index <= 6;
         when "1001010010100" => index <= 8;
         when "1001010010101" => index <= 7;
         when "1001010010110" => index <= 7;
         when "1001010010111" => index <= 6;
         when "1001010011000" => index <= 8;
         when "1001010011001" => index <= 7;
         when "1001010011010" => index <= 7;
         when "1001010011011" => index <= 6;
         when "1001010011100" => index <= 7;
         when "1001010011101" => index <= 6;
         when "1001010011110" => index <= 6;
         when "1001010011111" => index <= 6;
         when "1001010100000" => index <= 9;
         when "1001010100001" => index <= 8;
         when "1001010100010" => index <= 8;
         when "1001010100011" => index <= 7;
         when "1001010100100" => index <= 8;
         when "1001010100101" => index <= 7;
         when "1001010100110" => index <= 7;
         when "1001010100111" => index <= 6;
         when "1001010101000" => index <= 8;
         when "1001010101001" => index <= 7;
         when "1001010101010" => index <= 7;
         when "1001010101011" => index <= 6;
         when "1001010101100" => index <= 7;
         when "1001010101101" => index <= 6;
         when "1001010101110" => index <= 7;
         when "1001010101111" => index <= 6;
         when "1001010110000" => index <= 8;
         when "1001010110001" => index <= 7;
         when "1001010110010" => index <= 7;
         when "1001010110011" => index <= 6;
         when "1001010110100" => index <= 8;
         when "1001010110101" => index <= 7;
         when "1001010110110" => index <= 7;
         when "1001010110111" => index <= 6;
         when "1001010111000" => index <= 8;
         when "1001010111001" => index <= 7;
         when "1001010111010" => index <= 7;
         when "1001010111011" => index <= 6;
         when "1001010111100" => index <= 7;
         when "1001010111101" => index <= 6;
         when "1001010111110" => index <= 6;
         when "1001010111111" => index <= 6;
         when "1001011000000" => index <= 10;
         when "1001011000001" => index <= 8;
         when "1001011000010" => index <= 8;
         when "1001011000011" => index <= 7;
         when "1001011000100" => index <= 8;
         when "1001011000101" => index <= 7;
         when "1001011000110" => index <= 7;
         when "1001011000111" => index <= 6;
         when "1001011001000" => index <= 8;
         when "1001011001001" => index <= 7;
         when "1001011001010" => index <= 7;
         when "1001011001011" => index <= 6;
         when "1001011001100" => index <= 8;
         when "1001011001101" => index <= 7;
         when "1001011001110" => index <= 7;
         when "1001011001111" => index <= 6;
         when "1001011010000" => index <= 9;
         when "1001011010001" => index <= 7;
         when "1001011010010" => index <= 8;
         when "1001011010011" => index <= 7;
         when "1001011010100" => index <= 8;
         when "1001011010101" => index <= 7;
         when "1001011010110" => index <= 7;
         when "1001011010111" => index <= 6;
         when "1001011011000" => index <= 8;
         when "1001011011001" => index <= 7;
         when "1001011011010" => index <= 7;
         when "1001011011011" => index <= 6;
         when "1001011011100" => index <= 7;
         when "1001011011101" => index <= 6;
         when "1001011011110" => index <= 6;
         when "1001011011111" => index <= 6;
         when "1001011100000" => index <= 9;
         when "1001011100001" => index <= 8;
         when "1001011100010" => index <= 8;
         when "1001011100011" => index <= 7;
         when "1001011100100" => index <= 8;
         when "1001011100101" => index <= 7;
         when "1001011100110" => index <= 7;
         when "1001011100111" => index <= 6;
         when "1001011101000" => index <= 8;
         when "1001011101001" => index <= 7;
         when "1001011101010" => index <= 7;
         when "1001011101011" => index <= 6;
         when "1001011101100" => index <= 7;
         when "1001011101101" => index <= 6;
         when "1001011101110" => index <= 7;
         when "1001011101111" => index <= 6;
         when "1001011110000" => index <= 8;
         when "1001011110001" => index <= 7;
         when "1001011110010" => index <= 7;
         when "1001011110011" => index <= 6;
         when "1001011110100" => index <= 7;
         when "1001011110101" => index <= 7;
         when "1001011110110" => index <= 7;
         when "1001011110111" => index <= 6;
         when "1001011111000" => index <= 8;
         when "1001011111001" => index <= 7;
         when "1001011111010" => index <= 7;
         when "1001011111011" => index <= 6;
         when "1001011111100" => index <= 7;
         when "1001011111101" => index <= 6;
         when "1001011111110" => index <= 6;
         when "1001011111111" => index <= 6;
         when "1001100000000" => index <= 11;
         when "1001100000001" => index <= 8;
         when "1001100000010" => index <= 8;
         when "1001100000011" => index <= 7;
         when "1001100000100" => index <= 9;
         when "1001100000101" => index <= 7;
         when "1001100000110" => index <= 7;
         when "1001100000111" => index <= 6;
         when "1001100001000" => index <= 9;
         when "1001100001001" => index <= 7;
         when "1001100001010" => index <= 8;
         when "1001100001011" => index <= 6;
         when "1001100001100" => index <= 8;
         when "1001100001101" => index <= 7;
         when "1001100001110" => index <= 7;
         when "1001100001111" => index <= 6;
         when "1001100010000" => index <= 9;
         when "1001100010001" => index <= 8;
         when "1001100010010" => index <= 8;
         when "1001100010011" => index <= 7;
         when "1001100010100" => index <= 8;
         when "1001100010101" => index <= 7;
         when "1001100010110" => index <= 7;
         when "1001100010111" => index <= 6;
         when "1001100011000" => index <= 8;
         when "1001100011001" => index <= 7;
         when "1001100011010" => index <= 7;
         when "1001100011011" => index <= 6;
         when "1001100011100" => index <= 7;
         when "1001100011101" => index <= 6;
         when "1001100011110" => index <= 7;
         when "1001100011111" => index <= 6;
         when "1001100100000" => index <= 10;
         when "1001100100001" => index <= 8;
         when "1001100100010" => index <= 8;
         when "1001100100011" => index <= 7;
         when "1001100100100" => index <= 8;
         when "1001100100101" => index <= 7;
         when "1001100100110" => index <= 7;
         when "1001100100111" => index <= 6;
         when "1001100101000" => index <= 8;
         when "1001100101001" => index <= 7;
         when "1001100101010" => index <= 7;
         when "1001100101011" => index <= 6;
         when "1001100101100" => index <= 8;
         when "1001100101101" => index <= 7;
         when "1001100101110" => index <= 7;
         when "1001100101111" => index <= 6;
         when "1001100110000" => index <= 9;
         when "1001100110001" => index <= 7;
         when "1001100110010" => index <= 8;
         when "1001100110011" => index <= 7;
         when "1001100110100" => index <= 8;
         when "1001100110101" => index <= 7;
         when "1001100110110" => index <= 7;
         when "1001100110111" => index <= 6;
         when "1001100111000" => index <= 8;
         when "1001100111001" => index <= 7;
         when "1001100111010" => index <= 7;
         when "1001100111011" => index <= 6;
         when "1001100111100" => index <= 7;
         when "1001100111101" => index <= 6;
         when "1001100111110" => index <= 6;
         when "1001100111111" => index <= 6;
         when "1001101000000" => index <= 10;
         when "1001101000001" => index <= 8;
         when "1001101000010" => index <= 8;
         when "1001101000011" => index <= 7;
         when "1001101000100" => index <= 8;
         when "1001101000101" => index <= 7;
         when "1001101000110" => index <= 7;
         when "1001101000111" => index <= 6;
         when "1001101001000" => index <= 9;
         when "1001101001001" => index <= 7;
         when "1001101001010" => index <= 8;
         when "1001101001011" => index <= 7;
         when "1001101001100" => index <= 8;
         when "1001101001101" => index <= 7;
         when "1001101001110" => index <= 7;
         when "1001101001111" => index <= 6;
         when "1001101010000" => index <= 9;
         when "1001101010001" => index <= 8;
         when "1001101010010" => index <= 8;
         when "1001101010011" => index <= 7;
         when "1001101010100" => index <= 8;
         when "1001101010101" => index <= 7;
         when "1001101010110" => index <= 7;
         when "1001101010111" => index <= 6;
         when "1001101011000" => index <= 8;
         when "1001101011001" => index <= 7;
         when "1001101011010" => index <= 7;
         when "1001101011011" => index <= 6;
         when "1001101011100" => index <= 7;
         when "1001101011101" => index <= 6;
         when "1001101011110" => index <= 7;
         when "1001101011111" => index <= 6;
         when "1001101100000" => index <= 9;
         when "1001101100001" => index <= 8;
         when "1001101100010" => index <= 8;
         when "1001101100011" => index <= 7;
         when "1001101100100" => index <= 8;
         when "1001101100101" => index <= 7;
         when "1001101100110" => index <= 7;
         when "1001101100111" => index <= 6;
         when "1001101101000" => index <= 8;
         when "1001101101001" => index <= 7;
         when "1001101101010" => index <= 7;
         when "1001101101011" => index <= 6;
         when "1001101101100" => index <= 7;
         when "1001101101101" => index <= 7;
         when "1001101101110" => index <= 7;
         when "1001101101111" => index <= 6;
         when "1001101110000" => index <= 8;
         when "1001101110001" => index <= 7;
         when "1001101110010" => index <= 7;
         when "1001101110011" => index <= 7;
         when "1001101110100" => index <= 8;
         when "1001101110101" => index <= 7;
         when "1001101110110" => index <= 7;
         when "1001101110111" => index <= 6;
         when "1001101111000" => index <= 8;
         when "1001101111001" => index <= 7;
         when "1001101111010" => index <= 7;
         when "1001101111011" => index <= 6;
         when "1001101111100" => index <= 7;
         when "1001101111101" => index <= 6;
         when "1001101111110" => index <= 7;
         when "1001101111111" => index <= 6;
         when "1001110000000" => index <= 10;
         when "1001110000001" => index <= 8;
         when "1001110000010" => index <= 8;
         when "1001110000011" => index <= 7;
         when "1001110000100" => index <= 9;
         when "1001110000101" => index <= 7;
         when "1001110000110" => index <= 8;
         when "1001110000111" => index <= 7;
         when "1001110001000" => index <= 9;
         when "1001110001001" => index <= 8;
         when "1001110001010" => index <= 8;
         when "1001110001011" => index <= 7;
         when "1001110001100" => index <= 8;
         when "1001110001101" => index <= 7;
         when "1001110001110" => index <= 7;
         when "1001110001111" => index <= 6;
         when "1001110010000" => index <= 9;
         when "1001110010001" => index <= 8;
         when "1001110010010" => index <= 8;
         when "1001110010011" => index <= 7;
         when "1001110010100" => index <= 8;
         when "1001110010101" => index <= 7;
         when "1001110010110" => index <= 7;
         when "1001110010111" => index <= 6;
         when "1001110011000" => index <= 8;
         when "1001110011001" => index <= 7;
         when "1001110011010" => index <= 7;
         when "1001110011011" => index <= 6;
         when "1001110011100" => index <= 7;
         when "1001110011101" => index <= 7;
         when "1001110011110" => index <= 7;
         when "1001110011111" => index <= 6;
         when "1001110100000" => index <= 9;
         when "1001110100001" => index <= 8;
         when "1001110100010" => index <= 8;
         when "1001110100011" => index <= 7;
         when "1001110100100" => index <= 8;
         when "1001110100101" => index <= 7;
         when "1001110100110" => index <= 7;
         when "1001110100111" => index <= 6;
         when "1001110101000" => index <= 8;
         when "1001110101001" => index <= 7;
         when "1001110101010" => index <= 7;
         when "1001110101011" => index <= 7;
         when "1001110101100" => index <= 8;
         when "1001110101101" => index <= 7;
         when "1001110101110" => index <= 7;
         when "1001110101111" => index <= 6;
         when "1001110110000" => index <= 8;
         when "1001110110001" => index <= 7;
         when "1001110110010" => index <= 8;
         when "1001110110011" => index <= 7;
         when "1001110110100" => index <= 8;
         when "1001110110101" => index <= 7;
         when "1001110110110" => index <= 7;
         when "1001110110111" => index <= 6;
         when "1001110111000" => index <= 8;
         when "1001110111001" => index <= 7;
         when "1001110111010" => index <= 7;
         when "1001110111011" => index <= 6;
         when "1001110111100" => index <= 7;
         when "1001110111101" => index <= 7;
         when "1001110111110" => index <= 7;
         when "1001110111111" => index <= 6;
         when "1001111000000" => index <= 9;
         when "1001111000001" => index <= 8;
         when "1001111000010" => index <= 8;
         when "1001111000011" => index <= 7;
         when "1001111000100" => index <= 8;
         when "1001111000101" => index <= 7;
         when "1001111000110" => index <= 7;
         when "1001111000111" => index <= 7;
         when "1001111001000" => index <= 8;
         when "1001111001001" => index <= 7;
         when "1001111001010" => index <= 8;
         when "1001111001011" => index <= 7;
         when "1001111001100" => index <= 8;
         when "1001111001101" => index <= 7;
         when "1001111001110" => index <= 7;
         when "1001111001111" => index <= 6;
         when "1001111010000" => index <= 9;
         when "1001111010001" => index <= 8;
         when "1001111010010" => index <= 8;
         when "1001111010011" => index <= 7;
         when "1001111010100" => index <= 8;
         when "1001111010101" => index <= 7;
         when "1001111010110" => index <= 7;
         when "1001111010111" => index <= 6;
         when "1001111011000" => index <= 8;
         when "1001111011001" => index <= 7;
         when "1001111011010" => index <= 7;
         when "1001111011011" => index <= 7;
         when "1001111011100" => index <= 7;
         when "1001111011101" => index <= 7;
         when "1001111011110" => index <= 7;
         when "1001111011111" => index <= 6;
         when "1001111100000" => index <= 9;
         when "1001111100001" => index <= 8;
         when "1001111100010" => index <= 8;
         when "1001111100011" => index <= 7;
         when "1001111100100" => index <= 8;
         when "1001111100101" => index <= 7;
         when "1001111100110" => index <= 7;
         when "1001111100111" => index <= 7;
         when "1001111101000" => index <= 8;
         when "1001111101001" => index <= 7;
         when "1001111101010" => index <= 7;
         when "1001111101011" => index <= 7;
         when "1001111101100" => index <= 8;
         when "1001111101101" => index <= 7;
         when "1001111101110" => index <= 7;
         when "1001111101111" => index <= 6;
         when "1001111110000" => index <= 8;
         when "1001111110001" => index <= 7;
         when "1001111110010" => index <= 8;
         when "1001111110011" => index <= 7;
         when "1001111110100" => index <= 8;
         when "1001111110101" => index <= 7;
         when "1001111110110" => index <= 7;
         when "1001111110111" => index <= 6;
         when "1001111111000" => index <= 8;
         when "1001111111001" => index <= 7;
         when "1001111111010" => index <= 7;
         when "1001111111011" => index <= 6;
         when "1001111111100" => index <= 7;
         when "1001111111101" => index <= 7;
         when "1001111111110" => index <= 7;
         when "1001111111111" => index <= 6;
         when "1010000000000" => index <= 12;
         when "1010000000001" => index <= 8;
         when "1010000000010" => index <= 9;
         when "1010000000011" => index <= 7;
         when "1010000000100" => index <= 9;
         when "1010000000101" => index <= 7;
         when "1010000000110" => index <= 7;
         when "1010000000111" => index <= 6;
         when "1010000001000" => index <= 9;
         when "1010000001001" => index <= 7;
         when "1010000001010" => index <= 8;
         when "1010000001011" => index <= 6;
         when "1010000001100" => index <= 8;
         when "1010000001101" => index <= 6;
         when "1010000001110" => index <= 7;
         when "1010000001111" => index <= 6;
         when "1010000010000" => index <= 10;
         when "1010000010001" => index <= 8;
         when "1010000010010" => index <= 8;
         when "1010000010011" => index <= 6;
         when "1010000010100" => index <= 8;
         when "1010000010101" => index <= 7;
         when "1010000010110" => index <= 7;
         when "1010000010111" => index <= 6;
         when "1010000011000" => index <= 8;
         when "1010000011001" => index <= 7;
         when "1010000011010" => index <= 7;
         when "1010000011011" => index <= 6;
         when "1010000011100" => index <= 7;
         when "1010000011101" => index <= 6;
         when "1010000011110" => index <= 6;
         when "1010000011111" => index <= 6;
         when "1010000100000" => index <= 10;
         when "1010000100001" => index <= 8;
         when "1010000100010" => index <= 8;
         when "1010000100011" => index <= 7;
         when "1010000100100" => index <= 8;
         when "1010000100101" => index <= 7;
         when "1010000100110" => index <= 7;
         when "1010000100111" => index <= 6;
         when "1010000101000" => index <= 8;
         when "1010000101001" => index <= 7;
         when "1010000101010" => index <= 7;
         when "1010000101011" => index <= 6;
         when "1010000101100" => index <= 7;
         when "1010000101101" => index <= 6;
         when "1010000101110" => index <= 6;
         when "1010000101111" => index <= 6;
         when "1010000110000" => index <= 9;
         when "1010000110001" => index <= 7;
         when "1010000110010" => index <= 7;
         when "1010000110011" => index <= 6;
         when "1010000110100" => index <= 8;
         when "1010000110101" => index <= 6;
         when "1010000110110" => index <= 7;
         when "1010000110111" => index <= 6;
         when "1010000111000" => index <= 8;
         when "1010000111001" => index <= 7;
         when "1010000111010" => index <= 7;
         when "1010000111011" => index <= 6;
         when "1010000111100" => index <= 7;
         when "1010000111101" => index <= 6;
         when "1010000111110" => index <= 6;
         when "1010000111111" => index <= 6;
         when "1010001000000" => index <= 10;
         when "1010001000001" => index <= 8;
         when "1010001000010" => index <= 8;
         when "1010001000011" => index <= 7;
         when "1010001000100" => index <= 8;
         when "1010001000101" => index <= 7;
         when "1010001000110" => index <= 7;
         when "1010001000111" => index <= 6;
         when "1010001001000" => index <= 9;
         when "1010001001001" => index <= 7;
         when "1010001001010" => index <= 7;
         when "1010001001011" => index <= 6;
         when "1010001001100" => index <= 8;
         when "1010001001101" => index <= 6;
         when "1010001001110" => index <= 7;
         when "1010001001111" => index <= 6;
         when "1010001010000" => index <= 9;
         when "1010001010001" => index <= 7;
         when "1010001010010" => index <= 8;
         when "1010001010011" => index <= 6;
         when "1010001010100" => index <= 8;
         when "1010001010101" => index <= 7;
         when "1010001010110" => index <= 7;
         when "1010001010111" => index <= 6;
         when "1010001011000" => index <= 8;
         when "1010001011001" => index <= 7;
         when "1010001011010" => index <= 7;
         when "1010001011011" => index <= 6;
         when "1010001011100" => index <= 7;
         when "1010001011101" => index <= 6;
         when "1010001011110" => index <= 6;
         when "1010001011111" => index <= 6;
         when "1010001100000" => index <= 9;
         when "1010001100001" => index <= 8;
         when "1010001100010" => index <= 8;
         when "1010001100011" => index <= 7;
         when "1010001100100" => index <= 8;
         when "1010001100101" => index <= 7;
         when "1010001100110" => index <= 7;
         when "1010001100111" => index <= 6;
         when "1010001101000" => index <= 8;
         when "1010001101001" => index <= 7;
         when "1010001101010" => index <= 7;
         when "1010001101011" => index <= 6;
         when "1010001101100" => index <= 7;
         when "1010001101101" => index <= 6;
         when "1010001101110" => index <= 7;
         when "1010001101111" => index <= 6;
         when "1010001110000" => index <= 8;
         when "1010001110001" => index <= 7;
         when "1010001110010" => index <= 7;
         when "1010001110011" => index <= 6;
         when "1010001110100" => index <= 8;
         when "1010001110101" => index <= 7;
         when "1010001110110" => index <= 7;
         when "1010001110111" => index <= 6;
         when "1010001111000" => index <= 8;
         when "1010001111001" => index <= 7;
         when "1010001111010" => index <= 7;
         when "1010001111011" => index <= 6;
         when "1010001111100" => index <= 7;
         when "1010001111101" => index <= 6;
         when "1010001111110" => index <= 6;
         when "1010001111111" => index <= 6;
         when "1010010000000" => index <= 11;
         when "1010010000001" => index <= 8;
         when "1010010000010" => index <= 8;
         when "1010010000011" => index <= 7;
         when "1010010000100" => index <= 9;
         when "1010010000101" => index <= 7;
         when "1010010000110" => index <= 7;
         when "1010010000111" => index <= 6;
         when "1010010001000" => index <= 9;
         when "1010010001001" => index <= 7;
         when "1010010001010" => index <= 8;
         when "1010010001011" => index <= 6;
         when "1010010001100" => index <= 8;
         when "1010010001101" => index <= 7;
         when "1010010001110" => index <= 7;
         when "1010010001111" => index <= 6;
         when "1010010010000" => index <= 9;
         when "1010010010001" => index <= 8;
         when "1010010010010" => index <= 8;
         when "1010010010011" => index <= 7;
         when "1010010010100" => index <= 8;
         when "1010010010101" => index <= 7;
         when "1010010010110" => index <= 7;
         when "1010010010111" => index <= 6;
         when "1010010011000" => index <= 8;
         when "1010010011001" => index <= 7;
         when "1010010011010" => index <= 7;
         when "1010010011011" => index <= 6;
         when "1010010011100" => index <= 7;
         when "1010010011101" => index <= 6;
         when "1010010011110" => index <= 7;
         when "1010010011111" => index <= 6;
         when "1010010100000" => index <= 10;
         when "1010010100001" => index <= 8;
         when "1010010100010" => index <= 8;
         when "1010010100011" => index <= 7;
         when "1010010100100" => index <= 8;
         when "1010010100101" => index <= 7;
         when "1010010100110" => index <= 7;
         when "1010010100111" => index <= 6;
         when "1010010101000" => index <= 8;
         when "1010010101001" => index <= 7;
         when "1010010101010" => index <= 7;
         when "1010010101011" => index <= 6;
         when "1010010101100" => index <= 8;
         when "1010010101101" => index <= 7;
         when "1010010101110" => index <= 7;
         when "1010010101111" => index <= 6;
         when "1010010110000" => index <= 9;
         when "1010010110001" => index <= 7;
         when "1010010110010" => index <= 8;
         when "1010010110011" => index <= 7;
         when "1010010110100" => index <= 8;
         when "1010010110101" => index <= 7;
         when "1010010110110" => index <= 7;
         when "1010010110111" => index <= 6;
         when "1010010111000" => index <= 8;
         when "1010010111001" => index <= 7;
         when "1010010111010" => index <= 7;
         when "1010010111011" => index <= 6;
         when "1010010111100" => index <= 7;
         when "1010010111101" => index <= 6;
         when "1010010111110" => index <= 6;
         when "1010010111111" => index <= 6;
         when "1010011000000" => index <= 10;
         when "1010011000001" => index <= 8;
         when "1010011000010" => index <= 8;
         when "1010011000011" => index <= 7;
         when "1010011000100" => index <= 8;
         when "1010011000101" => index <= 7;
         when "1010011000110" => index <= 7;
         when "1010011000111" => index <= 6;
         when "1010011001000" => index <= 9;
         when "1010011001001" => index <= 7;
         when "1010011001010" => index <= 8;
         when "1010011001011" => index <= 7;
         when "1010011001100" => index <= 8;
         when "1010011001101" => index <= 7;
         when "1010011001110" => index <= 7;
         when "1010011001111" => index <= 6;
         when "1010011010000" => index <= 9;
         when "1010011010001" => index <= 8;
         when "1010011010010" => index <= 8;
         when "1010011010011" => index <= 7;
         when "1010011010100" => index <= 8;
         when "1010011010101" => index <= 7;
         when "1010011010110" => index <= 7;
         when "1010011010111" => index <= 6;
         when "1010011011000" => index <= 8;
         when "1010011011001" => index <= 7;
         when "1010011011010" => index <= 7;
         when "1010011011011" => index <= 6;
         when "1010011011100" => index <= 7;
         when "1010011011101" => index <= 6;
         when "1010011011110" => index <= 7;
         when "1010011011111" => index <= 6;
         when "1010011100000" => index <= 9;
         when "1010011100001" => index <= 8;
         when "1010011100010" => index <= 8;
         when "1010011100011" => index <= 7;
         when "1010011100100" => index <= 8;
         when "1010011100101" => index <= 7;
         when "1010011100110" => index <= 7;
         when "1010011100111" => index <= 6;
         when "1010011101000" => index <= 8;
         when "1010011101001" => index <= 7;
         when "1010011101010" => index <= 7;
         when "1010011101011" => index <= 6;
         when "1010011101100" => index <= 7;
         when "1010011101101" => index <= 7;
         when "1010011101110" => index <= 7;
         when "1010011101111" => index <= 6;
         when "1010011110000" => index <= 8;
         when "1010011110001" => index <= 7;
         when "1010011110010" => index <= 7;
         when "1010011110011" => index <= 7;
         when "1010011110100" => index <= 8;
         when "1010011110101" => index <= 7;
         when "1010011110110" => index <= 7;
         when "1010011110111" => index <= 6;
         when "1010011111000" => index <= 8;
         when "1010011111001" => index <= 7;
         when "1010011111010" => index <= 7;
         when "1010011111011" => index <= 6;
         when "1010011111100" => index <= 7;
         when "1010011111101" => index <= 6;
         when "1010011111110" => index <= 7;
         when "1010011111111" => index <= 6;
         when "1010100000000" => index <= 11;
         when "1010100000001" => index <= 8;
         when "1010100000010" => index <= 9;
         when "1010100000011" => index <= 7;
         when "1010100000100" => index <= 9;
         when "1010100000101" => index <= 7;
         when "1010100000110" => index <= 8;
         when "1010100000111" => index <= 6;
         when "1010100001000" => index <= 9;
         when "1010100001001" => index <= 8;
         when "1010100001010" => index <= 8;
         when "1010100001011" => index <= 7;
         when "1010100001100" => index <= 8;
         when "1010100001101" => index <= 7;
         when "1010100001110" => index <= 7;
         when "1010100001111" => index <= 6;
         when "1010100010000" => index <= 10;
         when "1010100010001" => index <= 8;
         when "1010100010010" => index <= 8;
         when "1010100010011" => index <= 7;
         when "1010100010100" => index <= 8;
         when "1010100010101" => index <= 7;
         when "1010100010110" => index <= 7;
         when "1010100010111" => index <= 6;
         when "1010100011000" => index <= 8;
         when "1010100011001" => index <= 7;
         when "1010100011010" => index <= 7;
         when "1010100011011" => index <= 6;
         when "1010100011100" => index <= 8;
         when "1010100011101" => index <= 7;
         when "1010100011110" => index <= 7;
         when "1010100011111" => index <= 6;
         when "1010100100000" => index <= 10;
         when "1010100100001" => index <= 8;
         when "1010100100010" => index <= 8;
         when "1010100100011" => index <= 7;
         when "1010100100100" => index <= 8;
         when "1010100100101" => index <= 7;
         when "1010100100110" => index <= 7;
         when "1010100100111" => index <= 6;
         when "1010100101000" => index <= 9;
         when "1010100101001" => index <= 7;
         when "1010100101010" => index <= 8;
         when "1010100101011" => index <= 7;
         when "1010100101100" => index <= 8;
         when "1010100101101" => index <= 7;
         when "1010100101110" => index <= 7;
         when "1010100101111" => index <= 6;
         when "1010100110000" => index <= 9;
         when "1010100110001" => index <= 8;
         when "1010100110010" => index <= 8;
         when "1010100110011" => index <= 7;
         when "1010100110100" => index <= 8;
         when "1010100110101" => index <= 7;
         when "1010100110110" => index <= 7;
         when "1010100110111" => index <= 6;
         when "1010100111000" => index <= 8;
         when "1010100111001" => index <= 7;
         when "1010100111010" => index <= 7;
         when "1010100111011" => index <= 6;
         when "1010100111100" => index <= 7;
         when "1010100111101" => index <= 6;
         when "1010100111110" => index <= 7;
         when "1010100111111" => index <= 6;
         when "1010101000000" => index <= 10;
         when "1010101000001" => index <= 8;
         when "1010101000010" => index <= 8;
         when "1010101000011" => index <= 7;
         when "1010101000100" => index <= 9;
         when "1010101000101" => index <= 7;
         when "1010101000110" => index <= 8;
         when "1010101000111" => index <= 7;
         when "1010101001000" => index <= 9;
         when "1010101001001" => index <= 8;
         when "1010101001010" => index <= 8;
         when "1010101001011" => index <= 7;
         when "1010101001100" => index <= 8;
         when "1010101001101" => index <= 7;
         when "1010101001110" => index <= 7;
         when "1010101001111" => index <= 6;
         when "1010101010000" => index <= 9;
         when "1010101010001" => index <= 8;
         when "1010101010010" => index <= 8;
         when "1010101010011" => index <= 7;
         when "1010101010100" => index <= 8;
         when "1010101010101" => index <= 7;
         when "1010101010110" => index <= 7;
         when "1010101010111" => index <= 6;
         when "1010101011000" => index <= 8;
         when "1010101011001" => index <= 7;
         when "1010101011010" => index <= 7;
         when "1010101011011" => index <= 6;
         when "1010101011100" => index <= 7;
         when "1010101011101" => index <= 7;
         when "1010101011110" => index <= 7;
         when "1010101011111" => index <= 6;
         when "1010101100000" => index <= 9;
         when "1010101100001" => index <= 8;
         when "1010101100010" => index <= 8;
         when "1010101100011" => index <= 7;
         when "1010101100100" => index <= 8;
         when "1010101100101" => index <= 7;
         when "1010101100110" => index <= 7;
         when "1010101100111" => index <= 6;
         when "1010101101000" => index <= 8;
         when "1010101101001" => index <= 7;
         when "1010101101010" => index <= 7;
         when "1010101101011" => index <= 7;
         when "1010101101100" => index <= 8;
         when "1010101101101" => index <= 7;
         when "1010101101110" => index <= 7;
         when "1010101101111" => index <= 6;
         when "1010101110000" => index <= 8;
         when "1010101110001" => index <= 7;
         when "1010101110010" => index <= 8;
         when "1010101110011" => index <= 7;
         when "1010101110100" => index <= 8;
         when "1010101110101" => index <= 7;
         when "1010101110110" => index <= 7;
         when "1010101110111" => index <= 6;
         when "1010101111000" => index <= 8;
         when "1010101111001" => index <= 7;
         when "1010101111010" => index <= 7;
         when "1010101111011" => index <= 6;
         when "1010101111100" => index <= 7;
         when "1010101111101" => index <= 7;
         when "1010101111110" => index <= 7;
         when "1010101111111" => index <= 6;
         when "1010110000000" => index <= 10;
         when "1010110000001" => index <= 8;
         when "1010110000010" => index <= 9;
         when "1010110000011" => index <= 7;
         when "1010110000100" => index <= 9;
         when "1010110000101" => index <= 8;
         when "1010110000110" => index <= 8;
         when "1010110000111" => index <= 7;
         when "1010110001000" => index <= 9;
         when "1010110001001" => index <= 8;
         when "1010110001010" => index <= 8;
         when "1010110001011" => index <= 7;
         when "1010110001100" => index <= 8;
         when "1010110001101" => index <= 7;
         when "1010110001110" => index <= 7;
         when "1010110001111" => index <= 6;
         when "1010110010000" => index <= 9;
         when "1010110010001" => index <= 8;
         when "1010110010010" => index <= 8;
         when "1010110010011" => index <= 7;
         when "1010110010100" => index <= 8;
         when "1010110010101" => index <= 7;
         when "1010110010110" => index <= 7;
         when "1010110010111" => index <= 6;
         when "1010110011000" => index <= 8;
         when "1010110011001" => index <= 7;
         when "1010110011010" => index <= 7;
         when "1010110011011" => index <= 7;
         when "1010110011100" => index <= 8;
         when "1010110011101" => index <= 7;
         when "1010110011110" => index <= 7;
         when "1010110011111" => index <= 6;
         when "1010110100000" => index <= 9;
         when "1010110100001" => index <= 8;
         when "1010110100010" => index <= 8;
         when "1010110100011" => index <= 7;
         when "1010110100100" => index <= 8;
         when "1010110100101" => index <= 7;
         when "1010110100110" => index <= 7;
         when "1010110100111" => index <= 7;
         when "1010110101000" => index <= 8;
         when "1010110101001" => index <= 7;
         when "1010110101010" => index <= 8;
         when "1010110101011" => index <= 7;
         when "1010110101100" => index <= 8;
         when "1010110101101" => index <= 7;
         when "1010110101110" => index <= 7;
         when "1010110101111" => index <= 6;
         when "1010110110000" => index <= 9;
         when "1010110110001" => index <= 8;
         when "1010110110010" => index <= 8;
         when "1010110110011" => index <= 7;
         when "1010110110100" => index <= 8;
         when "1010110110101" => index <= 7;
         when "1010110110110" => index <= 7;
         when "1010110110111" => index <= 6;
         when "1010110111000" => index <= 8;
         when "1010110111001" => index <= 7;
         when "1010110111010" => index <= 7;
         when "1010110111011" => index <= 7;
         when "1010110111100" => index <= 7;
         when "1010110111101" => index <= 7;
         when "1010110111110" => index <= 7;
         when "1010110111111" => index <= 6;
         when "1010111000000" => index <= 10;
         when "1010111000001" => index <= 8;
         when "1010111000010" => index <= 8;
         when "1010111000011" => index <= 7;
         when "1010111000100" => index <= 8;
         when "1010111000101" => index <= 7;
         when "1010111000110" => index <= 8;
         when "1010111000111" => index <= 7;
         when "1010111001000" => index <= 9;
         when "1010111001001" => index <= 8;
         when "1010111001010" => index <= 8;
         when "1010111001011" => index <= 7;
         when "1010111001100" => index <= 8;
         when "1010111001101" => index <= 7;
         when "1010111001110" => index <= 7;
         when "1010111001111" => index <= 6;
         when "1010111010000" => index <= 9;
         when "1010111010001" => index <= 8;
         when "1010111010010" => index <= 8;
         when "1010111010011" => index <= 7;
         when "1010111010100" => index <= 8;
         when "1010111010101" => index <= 7;
         when "1010111010110" => index <= 7;
         when "1010111010111" => index <= 7;
         when "1010111011000" => index <= 8;
         when "1010111011001" => index <= 7;
         when "1010111011010" => index <= 7;
         when "1010111011011" => index <= 7;
         when "1010111011100" => index <= 8;
         when "1010111011101" => index <= 7;
         when "1010111011110" => index <= 7;
         when "1010111011111" => index <= 6;
         when "1010111100000" => index <= 9;
         when "1010111100001" => index <= 8;
         when "1010111100010" => index <= 8;
         when "1010111100011" => index <= 7;
         when "1010111100100" => index <= 8;
         when "1010111100101" => index <= 7;
         when "1010111100110" => index <= 7;
         when "1010111100111" => index <= 7;
         when "1010111101000" => index <= 8;
         when "1010111101001" => index <= 7;
         when "1010111101010" => index <= 8;
         when "1010111101011" => index <= 7;
         when "1010111101100" => index <= 8;
         when "1010111101101" => index <= 7;
         when "1010111101110" => index <= 7;
         when "1010111101111" => index <= 6;
         when "1010111110000" => index <= 8;
         when "1010111110001" => index <= 8;
         when "1010111110010" => index <= 8;
         when "1010111110011" => index <= 7;
         when "1010111110100" => index <= 8;
         when "1010111110101" => index <= 7;
         when "1010111110110" => index <= 7;
         when "1010111110111" => index <= 6;
         when "1010111111000" => index <= 8;
         when "1010111111001" => index <= 7;
         when "1010111111010" => index <= 7;
         when "1010111111011" => index <= 7;
         when "1010111111100" => index <= 7;
         when "1010111111101" => index <= 7;
         when "1010111111110" => index <= 7;
         when "1010111111111" => index <= 6;
         when "1011000000000" => index <= 11;
         when "1011000000001" => index <= 9;
         when "1011000000010" => index <= 9;
         when "1011000000011" => index <= 7;
         when "1011000000100" => index <= 9;
         when "1011000000101" => index <= 8;
         when "1011000000110" => index <= 8;
         when "1011000000111" => index <= 7;
         when "1011000001000" => index <= 10;
         when "1011000001001" => index <= 8;
         when "1011000001010" => index <= 8;
         when "1011000001011" => index <= 7;
         when "1011000001100" => index <= 8;
         when "1011000001101" => index <= 7;
         when "1011000001110" => index <= 7;
         when "1011000001111" => index <= 6;
         when "1011000010000" => index <= 10;
         when "1011000010001" => index <= 8;
         when "1011000010010" => index <= 8;
         when "1011000010011" => index <= 7;
         when "1011000010100" => index <= 8;
         when "1011000010101" => index <= 7;
         when "1011000010110" => index <= 7;
         when "1011000010111" => index <= 6;
         when "1011000011000" => index <= 9;
         when "1011000011001" => index <= 7;
         when "1011000011010" => index <= 8;
         when "1011000011011" => index <= 7;
         when "1011000011100" => index <= 8;
         when "1011000011101" => index <= 7;
         when "1011000011110" => index <= 7;
         when "1011000011111" => index <= 6;
         when "1011000100000" => index <= 10;
         when "1011000100001" => index <= 8;
         when "1011000100010" => index <= 8;
         when "1011000100011" => index <= 7;
         when "1011000100100" => index <= 9;
         when "1011000100101" => index <= 7;
         when "1011000100110" => index <= 8;
         when "1011000100111" => index <= 7;
         when "1011000101000" => index <= 9;
         when "1011000101001" => index <= 8;
         when "1011000101010" => index <= 8;
         when "1011000101011" => index <= 7;
         when "1011000101100" => index <= 8;
         when "1011000101101" => index <= 7;
         when "1011000101110" => index <= 7;
         when "1011000101111" => index <= 6;
         when "1011000110000" => index <= 9;
         when "1011000110001" => index <= 8;
         when "1011000110010" => index <= 8;
         when "1011000110011" => index <= 7;
         when "1011000110100" => index <= 8;
         when "1011000110101" => index <= 7;
         when "1011000110110" => index <= 7;
         when "1011000110111" => index <= 6;
         when "1011000111000" => index <= 8;
         when "1011000111001" => index <= 7;
         when "1011000111010" => index <= 7;
         when "1011000111011" => index <= 6;
         when "1011000111100" => index <= 7;
         when "1011000111101" => index <= 7;
         when "1011000111110" => index <= 7;
         when "1011000111111" => index <= 6;
         when "1011001000000" => index <= 10;
         when "1011001000001" => index <= 8;
         when "1011001000010" => index <= 9;
         when "1011001000011" => index <= 7;
         when "1011001000100" => index <= 9;
         when "1011001000101" => index <= 8;
         when "1011001000110" => index <= 8;
         when "1011001000111" => index <= 7;
         when "1011001001000" => index <= 9;
         when "1011001001001" => index <= 8;
         when "1011001001010" => index <= 8;
         when "1011001001011" => index <= 7;
         when "1011001001100" => index <= 8;
         when "1011001001101" => index <= 7;
         when "1011001001110" => index <= 7;
         when "1011001001111" => index <= 6;
         when "1011001010000" => index <= 9;
         when "1011001010001" => index <= 8;
         when "1011001010010" => index <= 8;
         when "1011001010011" => index <= 7;
         when "1011001010100" => index <= 8;
         when "1011001010101" => index <= 7;
         when "1011001010110" => index <= 7;
         when "1011001010111" => index <= 6;
         when "1011001011000" => index <= 8;
         when "1011001011001" => index <= 7;
         when "1011001011010" => index <= 7;
         when "1011001011011" => index <= 7;
         when "1011001011100" => index <= 8;
         when "1011001011101" => index <= 7;
         when "1011001011110" => index <= 7;
         when "1011001011111" => index <= 6;
         when "1011001100000" => index <= 9;
         when "1011001100001" => index <= 8;
         when "1011001100010" => index <= 8;
         when "1011001100011" => index <= 7;
         when "1011001100100" => index <= 8;
         when "1011001100101" => index <= 7;
         when "1011001100110" => index <= 7;
         when "1011001100111" => index <= 7;
         when "1011001101000" => index <= 8;
         when "1011001101001" => index <= 7;
         when "1011001101010" => index <= 8;
         when "1011001101011" => index <= 7;
         when "1011001101100" => index <= 8;
         when "1011001101101" => index <= 7;
         when "1011001101110" => index <= 7;
         when "1011001101111" => index <= 6;
         when "1011001110000" => index <= 9;
         when "1011001110001" => index <= 8;
         when "1011001110010" => index <= 8;
         when "1011001110011" => index <= 7;
         when "1011001110100" => index <= 8;
         when "1011001110101" => index <= 7;
         when "1011001110110" => index <= 7;
         when "1011001110111" => index <= 6;
         when "1011001111000" => index <= 8;
         when "1011001111001" => index <= 7;
         when "1011001111010" => index <= 7;
         when "1011001111011" => index <= 7;
         when "1011001111100" => index <= 7;
         when "1011001111101" => index <= 7;
         when "1011001111110" => index <= 7;
         when "1011001111111" => index <= 6;
         when "1011010000000" => index <= 10;
         when "1011010000001" => index <= 9;
         when "1011010000010" => index <= 9;
         when "1011010000011" => index <= 8;
         when "1011010000100" => index <= 9;
         when "1011010000101" => index <= 8;
         when "1011010000110" => index <= 8;
         when "1011010000111" => index <= 7;
         when "1011010001000" => index <= 9;
         when "1011010001001" => index <= 8;
         when "1011010001010" => index <= 8;
         when "1011010001011" => index <= 7;
         when "1011010001100" => index <= 8;
         when "1011010001101" => index <= 7;
         when "1011010001110" => index <= 7;
         when "1011010001111" => index <= 6;
         when "1011010010000" => index <= 9;
         when "1011010010001" => index <= 8;
         when "1011010010010" => index <= 8;
         when "1011010010011" => index <= 7;
         when "1011010010100" => index <= 8;
         when "1011010010101" => index <= 7;
         when "1011010010110" => index <= 7;
         when "1011010010111" => index <= 7;
         when "1011010011000" => index <= 8;
         when "1011010011001" => index <= 7;
         when "1011010011010" => index <= 8;
         when "1011010011011" => index <= 7;
         when "1011010011100" => index <= 8;
         when "1011010011101" => index <= 7;
         when "1011010011110" => index <= 7;
         when "1011010011111" => index <= 6;
         when "1011010100000" => index <= 10;
         when "1011010100001" => index <= 8;
         when "1011010100010" => index <= 8;
         when "1011010100011" => index <= 7;
         when "1011010100100" => index <= 8;
         when "1011010100101" => index <= 7;
         when "1011010100110" => index <= 8;
         when "1011010100111" => index <= 7;
         when "1011010101000" => index <= 9;
         when "1011010101001" => index <= 8;
         when "1011010101010" => index <= 8;
         when "1011010101011" => index <= 7;
         when "1011010101100" => index <= 8;
         when "1011010101101" => index <= 7;
         when "1011010101110" => index <= 7;
         when "1011010101111" => index <= 6;
         when "1011010110000" => index <= 9;
         when "1011010110001" => index <= 8;
         when "1011010110010" => index <= 8;
         when "1011010110011" => index <= 7;
         when "1011010110100" => index <= 8;
         when "1011010110101" => index <= 7;
         when "1011010110110" => index <= 7;
         when "1011010110111" => index <= 7;
         when "1011010111000" => index <= 8;
         when "1011010111001" => index <= 7;
         when "1011010111010" => index <= 7;
         when "1011010111011" => index <= 7;
         when "1011010111100" => index <= 8;
         when "1011010111101" => index <= 7;
         when "1011010111110" => index <= 7;
         when "1011010111111" => index <= 6;
         when "1011011000000" => index <= 10;
         when "1011011000001" => index <= 8;
         when "1011011000010" => index <= 8;
         when "1011011000011" => index <= 7;
         when "1011011000100" => index <= 9;
         when "1011011000101" => index <= 8;
         when "1011011000110" => index <= 8;
         when "1011011000111" => index <= 7;
         when "1011011001000" => index <= 9;
         when "1011011001001" => index <= 8;
         when "1011011001010" => index <= 8;
         when "1011011001011" => index <= 7;
         when "1011011001100" => index <= 8;
         when "1011011001101" => index <= 7;
         when "1011011001110" => index <= 7;
         when "1011011001111" => index <= 7;
         when "1011011010000" => index <= 9;
         when "1011011010001" => index <= 8;
         when "1011011010010" => index <= 8;
         when "1011011010011" => index <= 7;
         when "1011011010100" => index <= 8;
         when "1011011010101" => index <= 7;
         when "1011011010110" => index <= 7;
         when "1011011010111" => index <= 7;
         when "1011011011000" => index <= 8;
         when "1011011011001" => index <= 7;
         when "1011011011010" => index <= 8;
         when "1011011011011" => index <= 7;
         when "1011011011100" => index <= 8;
         when "1011011011101" => index <= 7;
         when "1011011011110" => index <= 7;
         when "1011011011111" => index <= 6;
         when "1011011100000" => index <= 9;
         when "1011011100001" => index <= 8;
         when "1011011100010" => index <= 8;
         when "1011011100011" => index <= 7;
         when "1011011100100" => index <= 8;
         when "1011011100101" => index <= 7;
         when "1011011100110" => index <= 8;
         when "1011011100111" => index <= 7;
         when "1011011101000" => index <= 8;
         when "1011011101001" => index <= 8;
         when "1011011101010" => index <= 8;
         when "1011011101011" => index <= 7;
         when "1011011101100" => index <= 8;
         when "1011011101101" => index <= 7;
         when "1011011101110" => index <= 7;
         when "1011011101111" => index <= 6;
         when "1011011110000" => index <= 9;
         when "1011011110001" => index <= 8;
         when "1011011110010" => index <= 8;
         when "1011011110011" => index <= 7;
         when "1011011110100" => index <= 8;
         when "1011011110101" => index <= 7;
         when "1011011110110" => index <= 7;
         when "1011011110111" => index <= 7;
         when "1011011111000" => index <= 8;
         when "1011011111001" => index <= 7;
         when "1011011111010" => index <= 7;
         when "1011011111011" => index <= 7;
         when "1011011111100" => index <= 7;
         when "1011011111101" => index <= 7;
         when "1011011111110" => index <= 7;
         when "1011011111111" => index <= 6;
         when "1011100000000" => index <= 11;
         when "1011100000001" => index <= 9;
         when "1011100000010" => index <= 9;
         when "1011100000011" => index <= 8;
         when "1011100000100" => index <= 9;
         when "1011100000101" => index <= 8;
         when "1011100000110" => index <= 8;
         when "1011100000111" => index <= 7;
         when "1011100001000" => index <= 9;
         when "1011100001001" => index <= 8;
         when "1011100001010" => index <= 8;
         when "1011100001011" => index <= 7;
         when "1011100001100" => index <= 8;
         when "1011100001101" => index <= 7;
         when "1011100001110" => index <= 7;
         when "1011100001111" => index <= 7;
         when "1011100010000" => index <= 10;
         when "1011100010001" => index <= 8;
         when "1011100010010" => index <= 8;
         when "1011100010011" => index <= 7;
         when "1011100010100" => index <= 8;
         when "1011100010101" => index <= 7;
         when "1011100010110" => index <= 8;
         when "1011100010111" => index <= 7;
         when "1011100011000" => index <= 9;
         when "1011100011001" => index <= 8;
         when "1011100011010" => index <= 8;
         when "1011100011011" => index <= 7;
         when "1011100011100" => index <= 8;
         when "1011100011101" => index <= 7;
         when "1011100011110" => index <= 7;
         when "1011100011111" => index <= 6;
         when "1011100100000" => index <= 10;
         when "1011100100001" => index <= 8;
         when "1011100100010" => index <= 8;
         when "1011100100011" => index <= 7;
         when "1011100100100" => index <= 9;
         when "1011100100101" => index <= 8;
         when "1011100100110" => index <= 8;
         when "1011100100111" => index <= 7;
         when "1011100101000" => index <= 9;
         when "1011100101001" => index <= 8;
         when "1011100101010" => index <= 8;
         when "1011100101011" => index <= 7;
         when "1011100101100" => index <= 8;
         when "1011100101101" => index <= 7;
         when "1011100101110" => index <= 7;
         when "1011100101111" => index <= 7;
         when "1011100110000" => index <= 9;
         when "1011100110001" => index <= 8;
         when "1011100110010" => index <= 8;
         when "1011100110011" => index <= 7;
         when "1011100110100" => index <= 8;
         when "1011100110101" => index <= 7;
         when "1011100110110" => index <= 7;
         when "1011100110111" => index <= 7;
         when "1011100111000" => index <= 8;
         when "1011100111001" => index <= 7;
         when "1011100111010" => index <= 8;
         when "1011100111011" => index <= 7;
         when "1011100111100" => index <= 8;
         when "1011100111101" => index <= 7;
         when "1011100111110" => index <= 7;
         when "1011100111111" => index <= 6;
         when "1011101000000" => index <= 10;
         when "1011101000001" => index <= 8;
         when "1011101000010" => index <= 9;
         when "1011101000011" => index <= 8;
         when "1011101000100" => index <= 9;
         when "1011101000101" => index <= 8;
         when "1011101000110" => index <= 8;
         when "1011101000111" => index <= 7;
         when "1011101001000" => index <= 9;
         when "1011101001001" => index <= 8;
         when "1011101001010" => index <= 8;
         when "1011101001011" => index <= 7;
         when "1011101001100" => index <= 8;
         when "1011101001101" => index <= 7;
         when "1011101001110" => index <= 7;
         when "1011101001111" => index <= 7;
         when "1011101010000" => index <= 9;
         when "1011101010001" => index <= 8;
         when "1011101010010" => index <= 8;
         when "1011101010011" => index <= 7;
         when "1011101010100" => index <= 8;
         when "1011101010101" => index <= 7;
         when "1011101010110" => index <= 8;
         when "1011101010111" => index <= 7;
         when "1011101011000" => index <= 8;
         when "1011101011001" => index <= 8;
         when "1011101011010" => index <= 8;
         when "1011101011011" => index <= 7;
         when "1011101011100" => index <= 8;
         when "1011101011101" => index <= 7;
         when "1011101011110" => index <= 7;
         when "1011101011111" => index <= 6;
         when "1011101100000" => index <= 9;
         when "1011101100001" => index <= 8;
         when "1011101100010" => index <= 8;
         when "1011101100011" => index <= 7;
         when "1011101100100" => index <= 8;
         when "1011101100101" => index <= 8;
         when "1011101100110" => index <= 8;
         when "1011101100111" => index <= 7;
         when "1011101101000" => index <= 9;
         when "1011101101001" => index <= 8;
         when "1011101101010" => index <= 8;
         when "1011101101011" => index <= 7;
         when "1011101101100" => index <= 8;
         when "1011101101101" => index <= 7;
         when "1011101101110" => index <= 7;
         when "1011101101111" => index <= 7;
         when "1011101110000" => index <= 9;
         when "1011101110001" => index <= 8;
         when "1011101110010" => index <= 8;
         when "1011101110011" => index <= 7;
         when "1011101110100" => index <= 8;
         when "1011101110101" => index <= 7;
         when "1011101110110" => index <= 7;
         when "1011101110111" => index <= 7;
         when "1011101111000" => index <= 8;
         when "1011101111001" => index <= 7;
         when "1011101111010" => index <= 7;
         when "1011101111011" => index <= 7;
         when "1011101111100" => index <= 8;
         when "1011101111101" => index <= 7;
         when "1011101111110" => index <= 7;
         when "1011101111111" => index <= 6;
         when "1011110000000" => index <= 10;
         when "1011110000001" => index <= 9;
         when "1011110000010" => index <= 9;
         when "1011110000011" => index <= 8;
         when "1011110000100" => index <= 9;
         when "1011110000101" => index <= 8;
         when "1011110000110" => index <= 8;
         when "1011110000111" => index <= 7;
         when "1011110001000" => index <= 9;
         when "1011110001001" => index <= 8;
         when "1011110001010" => index <= 8;
         when "1011110001011" => index <= 7;
         when "1011110001100" => index <= 8;
         when "1011110001101" => index <= 7;
         when "1011110001110" => index <= 8;
         when "1011110001111" => index <= 7;
         when "1011110010000" => index <= 9;
         when "1011110010001" => index <= 8;
         when "1011110010010" => index <= 8;
         when "1011110010011" => index <= 7;
         when "1011110010100" => index <= 8;
         when "1011110010101" => index <= 8;
         when "1011110010110" => index <= 8;
         when "1011110010111" => index <= 7;
         when "1011110011000" => index <= 9;
         when "1011110011001" => index <= 8;
         when "1011110011010" => index <= 8;
         when "1011110011011" => index <= 7;
         when "1011110011100" => index <= 8;
         when "1011110011101" => index <= 7;
         when "1011110011110" => index <= 7;
         when "1011110011111" => index <= 7;
         when "1011110100000" => index <= 10;
         when "1011110100001" => index <= 8;
         when "1011110100010" => index <= 8;
         when "1011110100011" => index <= 8;
         when "1011110100100" => index <= 9;
         when "1011110100101" => index <= 8;
         when "1011110100110" => index <= 8;
         when "1011110100111" => index <= 7;
         when "1011110101000" => index <= 9;
         when "1011110101001" => index <= 8;
         when "1011110101010" => index <= 8;
         when "1011110101011" => index <= 7;
         when "1011110101100" => index <= 8;
         when "1011110101101" => index <= 7;
         when "1011110101110" => index <= 7;
         when "1011110101111" => index <= 7;
         when "1011110110000" => index <= 9;
         when "1011110110001" => index <= 8;
         when "1011110110010" => index <= 8;
         when "1011110110011" => index <= 7;
         when "1011110110100" => index <= 8;
         when "1011110110101" => index <= 7;
         when "1011110110110" => index <= 7;
         when "1011110110111" => index <= 7;
         when "1011110111000" => index <= 8;
         when "1011110111001" => index <= 7;
         when "1011110111010" => index <= 8;
         when "1011110111011" => index <= 7;
         when "1011110111100" => index <= 8;
         when "1011110111101" => index <= 7;
         when "1011110111110" => index <= 7;
         when "1011110111111" => index <= 7;
         when "1011111000000" => index <= 10;
         when "1011111000001" => index <= 8;
         when "1011111000010" => index <= 9;
         when "1011111000011" => index <= 8;
         when "1011111000100" => index <= 9;
         when "1011111000101" => index <= 8;
         when "1011111000110" => index <= 8;
         when "1011111000111" => index <= 7;
         when "1011111001000" => index <= 9;
         when "1011111001001" => index <= 8;
         when "1011111001010" => index <= 8;
         when "1011111001011" => index <= 7;
         when "1011111001100" => index <= 8;
         when "1011111001101" => index <= 7;
         when "1011111001110" => index <= 7;
         when "1011111001111" => index <= 7;
         when "1011111010000" => index <= 9;
         when "1011111010001" => index <= 8;
         when "1011111010010" => index <= 8;
         when "1011111010011" => index <= 7;
         when "1011111010100" => index <= 8;
         when "1011111010101" => index <= 7;
         when "1011111010110" => index <= 8;
         when "1011111010111" => index <= 7;
         when "1011111011000" => index <= 8;
         when "1011111011001" => index <= 8;
         when "1011111011010" => index <= 8;
         when "1011111011011" => index <= 7;
         when "1011111011100" => index <= 8;
         when "1011111011101" => index <= 7;
         when "1011111011110" => index <= 7;
         when "1011111011111" => index <= 7;
         when "1011111100000" => index <= 9;
         when "1011111100001" => index <= 8;
         when "1011111100010" => index <= 8;
         when "1011111100011" => index <= 7;
         when "1011111100100" => index <= 8;
         when "1011111100101" => index <= 8;
         when "1011111100110" => index <= 8;
         when "1011111100111" => index <= 7;
         when "1011111101000" => index <= 8;
         when "1011111101001" => index <= 8;
         when "1011111101010" => index <= 8;
         when "1011111101011" => index <= 7;
         when "1011111101100" => index <= 8;
         when "1011111101101" => index <= 7;
         when "1011111101110" => index <= 7;
         when "1011111101111" => index <= 7;
         when "1011111110000" => index <= 9;
         when "1011111110001" => index <= 8;
         when "1011111110010" => index <= 8;
         when "1011111110011" => index <= 7;
         when "1011111110100" => index <= 8;
         when "1011111110101" => index <= 7;
         when "1011111110110" => index <= 7;
         when "1011111110111" => index <= 7;
         when "1011111111000" => index <= 8;
         when "1011111111001" => index <= 7;
         when "1011111111010" => index <= 8;
         when "1011111111011" => index <= 7;
         when "1011111111100" => index <= 8;
         when "1011111111101" => index <= 7;
         when "1011111111110" => index <= 7;
         when "1011111111111" => index <= 7;
         when "1100000000000" => index <= 12;
         when "1100000000001" => index <= 9;
         when "1100000000010" => index <= 9;
         when "1100000000011" => index <= 7;
         when "1100000000100" => index <= 9;
         when "1100000000101" => index <= 7;
         when "1100000000110" => index <= 8;
         when "1100000000111" => index <= 6;
         when "1100000001000" => index <= 10;
         when "1100000001001" => index <= 8;
         when "1100000001010" => index <= 8;
         when "1100000001011" => index <= 6;
         when "1100000001100" => index <= 8;
         when "1100000001101" => index <= 7;
         when "1100000001110" => index <= 7;
         when "1100000001111" => index <= 6;
         when "1100000010000" => index <= 10;
         when "1100000010001" => index <= 8;
         when "1100000010010" => index <= 8;
         when "1100000010011" => index <= 7;
         when "1100000010100" => index <= 8;
         when "1100000010101" => index <= 7;
         when "1100000010110" => index <= 7;
         when "1100000010111" => index <= 6;
         when "1100000011000" => index <= 8;
         when "1100000011001" => index <= 7;
         when "1100000011010" => index <= 7;
         when "1100000011011" => index <= 6;
         when "1100000011100" => index <= 7;
         when "1100000011101" => index <= 6;
         when "1100000011110" => index <= 6;
         when "1100000011111" => index <= 6;
         when "1100000100000" => index <= 10;
         when "1100000100001" => index <= 8;
         when "1100000100010" => index <= 8;
         when "1100000100011" => index <= 7;
         when "1100000100100" => index <= 8;
         when "1100000100101" => index <= 7;
         when "1100000100110" => index <= 7;
         when "1100000100111" => index <= 6;
         when "1100000101000" => index <= 9;
         when "1100000101001" => index <= 7;
         when "1100000101010" => index <= 7;
         when "1100000101011" => index <= 6;
         when "1100000101100" => index <= 8;
         when "1100000101101" => index <= 6;
         when "1100000101110" => index <= 7;
         when "1100000101111" => index <= 6;
         when "1100000110000" => index <= 9;
         when "1100000110001" => index <= 7;
         when "1100000110010" => index <= 8;
         when "1100000110011" => index <= 6;
         when "1100000110100" => index <= 8;
         when "1100000110101" => index <= 7;
         when "1100000110110" => index <= 7;
         when "1100000110111" => index <= 6;
         when "1100000111000" => index <= 8;
         when "1100000111001" => index <= 7;
         when "1100000111010" => index <= 7;
         when "1100000111011" => index <= 6;
         when "1100000111100" => index <= 7;
         when "1100000111101" => index <= 6;
         when "1100000111110" => index <= 6;
         when "1100000111111" => index <= 6;
         when "1100001000000" => index <= 11;
         when "1100001000001" => index <= 8;
         when "1100001000010" => index <= 8;
         when "1100001000011" => index <= 7;
         when "1100001000100" => index <= 9;
         when "1100001000101" => index <= 7;
         when "1100001000110" => index <= 7;
         when "1100001000111" => index <= 6;
         when "1100001001000" => index <= 9;
         when "1100001001001" => index <= 7;
         when "1100001001010" => index <= 8;
         when "1100001001011" => index <= 6;
         when "1100001001100" => index <= 8;
         when "1100001001101" => index <= 7;
         when "1100001001110" => index <= 7;
         when "1100001001111" => index <= 6;
         when "1100001010000" => index <= 9;
         when "1100001010001" => index <= 8;
         when "1100001010010" => index <= 8;
         when "1100001010011" => index <= 7;
         when "1100001010100" => index <= 8;
         when "1100001010101" => index <= 7;
         when "1100001010110" => index <= 7;
         when "1100001010111" => index <= 6;
         when "1100001011000" => index <= 8;
         when "1100001011001" => index <= 7;
         when "1100001011010" => index <= 7;
         when "1100001011011" => index <= 6;
         when "1100001011100" => index <= 7;
         when "1100001011101" => index <= 6;
         when "1100001011110" => index <= 7;
         when "1100001011111" => index <= 6;
         when "1100001100000" => index <= 10;
         when "1100001100001" => index <= 8;
         when "1100001100010" => index <= 8;
         when "1100001100011" => index <= 7;
         when "1100001100100" => index <= 8;
         when "1100001100101" => index <= 7;
         when "1100001100110" => index <= 7;
         when "1100001100111" => index <= 6;
         when "1100001101000" => index <= 8;
         when "1100001101001" => index <= 7;
         when "1100001101010" => index <= 7;
         when "1100001101011" => index <= 6;
         when "1100001101100" => index <= 8;
         when "1100001101101" => index <= 7;
         when "1100001101110" => index <= 7;
         when "1100001101111" => index <= 6;
         when "1100001110000" => index <= 9;
         when "1100001110001" => index <= 7;
         when "1100001110010" => index <= 8;
         when "1100001110011" => index <= 7;
         when "1100001110100" => index <= 8;
         when "1100001110101" => index <= 7;
         when "1100001110110" => index <= 7;
         when "1100001110111" => index <= 6;
         when "1100001111000" => index <= 8;
         when "1100001111001" => index <= 7;
         when "1100001111010" => index <= 7;
         when "1100001111011" => index <= 6;
         when "1100001111100" => index <= 7;
         when "1100001111101" => index <= 6;
         when "1100001111110" => index <= 6;
         when "1100001111111" => index <= 6;
         when "1100010000000" => index <= 11;
         when "1100010000001" => index <= 8;
         when "1100010000010" => index <= 9;
         when "1100010000011" => index <= 7;
         when "1100010000100" => index <= 9;
         when "1100010000101" => index <= 7;
         when "1100010000110" => index <= 8;
         when "1100010000111" => index <= 6;
         when "1100010001000" => index <= 9;
         when "1100010001001" => index <= 8;
         when "1100010001010" => index <= 8;
         when "1100010001011" => index <= 7;
         when "1100010001100" => index <= 8;
         when "1100010001101" => index <= 7;
         when "1100010001110" => index <= 7;
         when "1100010001111" => index <= 6;
         when "1100010010000" => index <= 10;
         when "1100010010001" => index <= 8;
         when "1100010010010" => index <= 8;
         when "1100010010011" => index <= 7;
         when "1100010010100" => index <= 8;
         when "1100010010101" => index <= 7;
         when "1100010010110" => index <= 7;
         when "1100010010111" => index <= 6;
         when "1100010011000" => index <= 8;
         when "1100010011001" => index <= 7;
         when "1100010011010" => index <= 7;
         when "1100010011011" => index <= 6;
         when "1100010011100" => index <= 8;
         when "1100010011101" => index <= 7;
         when "1100010011110" => index <= 7;
         when "1100010011111" => index <= 6;
         when "1100010100000" => index <= 10;
         when "1100010100001" => index <= 8;
         when "1100010100010" => index <= 8;
         when "1100010100011" => index <= 7;
         when "1100010100100" => index <= 8;
         when "1100010100101" => index <= 7;
         when "1100010100110" => index <= 7;
         when "1100010100111" => index <= 6;
         when "1100010101000" => index <= 9;
         when "1100010101001" => index <= 7;
         when "1100010101010" => index <= 8;
         when "1100010101011" => index <= 7;
         when "1100010101100" => index <= 8;
         when "1100010101101" => index <= 7;
         when "1100010101110" => index <= 7;
         when "1100010101111" => index <= 6;
         when "1100010110000" => index <= 9;
         when "1100010110001" => index <= 8;
         when "1100010110010" => index <= 8;
         when "1100010110011" => index <= 7;
         when "1100010110100" => index <= 8;
         when "1100010110101" => index <= 7;
         when "1100010110110" => index <= 7;
         when "1100010110111" => index <= 6;
         when "1100010111000" => index <= 8;
         when "1100010111001" => index <= 7;
         when "1100010111010" => index <= 7;
         when "1100010111011" => index <= 6;
         when "1100010111100" => index <= 7;
         when "1100010111101" => index <= 6;
         when "1100010111110" => index <= 7;
         when "1100010111111" => index <= 6;
         when "1100011000000" => index <= 10;
         when "1100011000001" => index <= 8;
         when "1100011000010" => index <= 8;
         when "1100011000011" => index <= 7;
         when "1100011000100" => index <= 9;
         when "1100011000101" => index <= 7;
         when "1100011000110" => index <= 8;
         when "1100011000111" => index <= 7;
         when "1100011001000" => index <= 9;
         when "1100011001001" => index <= 8;
         when "1100011001010" => index <= 8;
         when "1100011001011" => index <= 7;
         when "1100011001100" => index <= 8;
         when "1100011001101" => index <= 7;
         when "1100011001110" => index <= 7;
         when "1100011001111" => index <= 6;
         when "1100011010000" => index <= 9;
         when "1100011010001" => index <= 8;
         when "1100011010010" => index <= 8;
         when "1100011010011" => index <= 7;
         when "1100011010100" => index <= 8;
         when "1100011010101" => index <= 7;
         when "1100011010110" => index <= 7;
         when "1100011010111" => index <= 6;
         when "1100011011000" => index <= 8;
         when "1100011011001" => index <= 7;
         when "1100011011010" => index <= 7;
         when "1100011011011" => index <= 6;
         when "1100011011100" => index <= 7;
         when "1100011011101" => index <= 7;
         when "1100011011110" => index <= 7;
         when "1100011011111" => index <= 6;
         when "1100011100000" => index <= 9;
         when "1100011100001" => index <= 8;
         when "1100011100010" => index <= 8;
         when "1100011100011" => index <= 7;
         when "1100011100100" => index <= 8;
         when "1100011100101" => index <= 7;
         when "1100011100110" => index <= 7;
         when "1100011100111" => index <= 6;
         when "1100011101000" => index <= 8;
         when "1100011101001" => index <= 7;
         when "1100011101010" => index <= 7;
         when "1100011101011" => index <= 7;
         when "1100011101100" => index <= 8;
         when "1100011101101" => index <= 7;
         when "1100011101110" => index <= 7;
         when "1100011101111" => index <= 6;
         when "1100011110000" => index <= 8;
         when "1100011110001" => index <= 7;
         when "1100011110010" => index <= 8;
         when "1100011110011" => index <= 7;
         when "1100011110100" => index <= 8;
         when "1100011110101" => index <= 7;
         when "1100011110110" => index <= 7;
         when "1100011110111" => index <= 6;
         when "1100011111000" => index <= 8;
         when "1100011111001" => index <= 7;
         when "1100011111010" => index <= 7;
         when "1100011111011" => index <= 6;
         when "1100011111100" => index <= 7;
         when "1100011111101" => index <= 7;
         when "1100011111110" => index <= 7;
         when "1100011111111" => index <= 6;
         when "1100100000000" => index <= 11;
         when "1100100000001" => index <= 9;
         when "1100100000010" => index <= 9;
         when "1100100000011" => index <= 7;
         when "1100100000100" => index <= 9;
         when "1100100000101" => index <= 8;
         when "1100100000110" => index <= 8;
         when "1100100000111" => index <= 7;
         when "1100100001000" => index <= 10;
         when "1100100001001" => index <= 8;
         when "1100100001010" => index <= 8;
         when "1100100001011" => index <= 7;
         when "1100100001100" => index <= 8;
         when "1100100001101" => index <= 7;
         when "1100100001110" => index <= 7;
         when "1100100001111" => index <= 6;
         when "1100100010000" => index <= 10;
         when "1100100010001" => index <= 8;
         when "1100100010010" => index <= 8;
         when "1100100010011" => index <= 7;
         when "1100100010100" => index <= 8;
         when "1100100010101" => index <= 7;
         when "1100100010110" => index <= 7;
         when "1100100010111" => index <= 6;
         when "1100100011000" => index <= 9;
         when "1100100011001" => index <= 7;
         when "1100100011010" => index <= 8;
         when "1100100011011" => index <= 7;
         when "1100100011100" => index <= 8;
         when "1100100011101" => index <= 7;
         when "1100100011110" => index <= 7;
         when "1100100011111" => index <= 6;
         when "1100100100000" => index <= 10;
         when "1100100100001" => index <= 8;
         when "1100100100010" => index <= 8;
         when "1100100100011" => index <= 7;
         when "1100100100100" => index <= 9;
         when "1100100100101" => index <= 7;
         when "1100100100110" => index <= 8;
         when "1100100100111" => index <= 7;
         when "1100100101000" => index <= 9;
         when "1100100101001" => index <= 8;
         when "1100100101010" => index <= 8;
         when "1100100101011" => index <= 7;
         when "1100100101100" => index <= 8;
         when "1100100101101" => index <= 7;
         when "1100100101110" => index <= 7;
         when "1100100101111" => index <= 6;
         when "1100100110000" => index <= 9;
         when "1100100110001" => index <= 8;
         when "1100100110010" => index <= 8;
         when "1100100110011" => index <= 7;
         when "1100100110100" => index <= 8;
         when "1100100110101" => index <= 7;
         when "1100100110110" => index <= 7;
         when "1100100110111" => index <= 6;
         when "1100100111000" => index <= 8;
         when "1100100111001" => index <= 7;
         when "1100100111010" => index <= 7;
         when "1100100111011" => index <= 6;
         when "1100100111100" => index <= 7;
         when "1100100111101" => index <= 7;
         when "1100100111110" => index <= 7;
         when "1100100111111" => index <= 6;
         when "1100101000000" => index <= 10;
         when "1100101000001" => index <= 8;
         when "1100101000010" => index <= 9;
         when "1100101000011" => index <= 7;
         when "1100101000100" => index <= 9;
         when "1100101000101" => index <= 8;
         when "1100101000110" => index <= 8;
         when "1100101000111" => index <= 7;
         when "1100101001000" => index <= 9;
         when "1100101001001" => index <= 8;
         when "1100101001010" => index <= 8;
         when "1100101001011" => index <= 7;
         when "1100101001100" => index <= 8;
         when "1100101001101" => index <= 7;
         when "1100101001110" => index <= 7;
         when "1100101001111" => index <= 6;
         when "1100101010000" => index <= 9;
         when "1100101010001" => index <= 8;
         when "1100101010010" => index <= 8;
         when "1100101010011" => index <= 7;
         when "1100101010100" => index <= 8;
         when "1100101010101" => index <= 7;
         when "1100101010110" => index <= 7;
         when "1100101010111" => index <= 6;
         when "1100101011000" => index <= 8;
         when "1100101011001" => index <= 7;
         when "1100101011010" => index <= 7;
         when "1100101011011" => index <= 7;
         when "1100101011100" => index <= 8;
         when "1100101011101" => index <= 7;
         when "1100101011110" => index <= 7;
         when "1100101011111" => index <= 6;
         when "1100101100000" => index <= 9;
         when "1100101100001" => index <= 8;
         when "1100101100010" => index <= 8;
         when "1100101100011" => index <= 7;
         when "1100101100100" => index <= 8;
         when "1100101100101" => index <= 7;
         when "1100101100110" => index <= 7;
         when "1100101100111" => index <= 7;
         when "1100101101000" => index <= 8;
         when "1100101101001" => index <= 7;
         when "1100101101010" => index <= 8;
         when "1100101101011" => index <= 7;
         when "1100101101100" => index <= 8;
         when "1100101101101" => index <= 7;
         when "1100101101110" => index <= 7;
         when "1100101101111" => index <= 6;
         when "1100101110000" => index <= 9;
         when "1100101110001" => index <= 8;
         when "1100101110010" => index <= 8;
         when "1100101110011" => index <= 7;
         when "1100101110100" => index <= 8;
         when "1100101110101" => index <= 7;
         when "1100101110110" => index <= 7;
         when "1100101110111" => index <= 6;
         when "1100101111000" => index <= 8;
         when "1100101111001" => index <= 7;
         when "1100101111010" => index <= 7;
         when "1100101111011" => index <= 7;
         when "1100101111100" => index <= 7;
         when "1100101111101" => index <= 7;
         when "1100101111110" => index <= 7;
         when "1100101111111" => index <= 6;
         when "1100110000000" => index <= 10;
         when "1100110000001" => index <= 9;
         when "1100110000010" => index <= 9;
         when "1100110000011" => index <= 8;
         when "1100110000100" => index <= 9;
         when "1100110000101" => index <= 8;
         when "1100110000110" => index <= 8;
         when "1100110000111" => index <= 7;
         when "1100110001000" => index <= 9;
         when "1100110001001" => index <= 8;
         when "1100110001010" => index <= 8;
         when "1100110001011" => index <= 7;
         when "1100110001100" => index <= 8;
         when "1100110001101" => index <= 7;
         when "1100110001110" => index <= 7;
         when "1100110001111" => index <= 6;
         when "1100110010000" => index <= 9;
         when "1100110010001" => index <= 8;
         when "1100110010010" => index <= 8;
         when "1100110010011" => index <= 7;
         when "1100110010100" => index <= 8;
         when "1100110010101" => index <= 7;
         when "1100110010110" => index <= 7;
         when "1100110010111" => index <= 7;
         when "1100110011000" => index <= 8;
         when "1100110011001" => index <= 7;
         when "1100110011010" => index <= 8;
         when "1100110011011" => index <= 7;
         when "1100110011100" => index <= 8;
         when "1100110011101" => index <= 7;
         when "1100110011110" => index <= 7;
         when "1100110011111" => index <= 6;
         when "1100110100000" => index <= 10;
         when "1100110100001" => index <= 8;
         when "1100110100010" => index <= 8;
         when "1100110100011" => index <= 7;
         when "1100110100100" => index <= 8;
         when "1100110100101" => index <= 7;
         when "1100110100110" => index <= 8;
         when "1100110100111" => index <= 7;
         when "1100110101000" => index <= 9;
         when "1100110101001" => index <= 8;
         when "1100110101010" => index <= 8;
         when "1100110101011" => index <= 7;
         when "1100110101100" => index <= 8;
         when "1100110101101" => index <= 7;
         when "1100110101110" => index <= 7;
         when "1100110101111" => index <= 6;
         when "1100110110000" => index <= 9;
         when "1100110110001" => index <= 8;
         when "1100110110010" => index <= 8;
         when "1100110110011" => index <= 7;
         when "1100110110100" => index <= 8;
         when "1100110110101" => index <= 7;
         when "1100110110110" => index <= 7;
         when "1100110110111" => index <= 7;
         when "1100110111000" => index <= 8;
         when "1100110111001" => index <= 7;
         when "1100110111010" => index <= 7;
         when "1100110111011" => index <= 7;
         when "1100110111100" => index <= 8;
         when "1100110111101" => index <= 7;
         when "1100110111110" => index <= 7;
         when "1100110111111" => index <= 6;
         when "1100111000000" => index <= 10;
         when "1100111000001" => index <= 8;
         when "1100111000010" => index <= 8;
         when "1100111000011" => index <= 7;
         when "1100111000100" => index <= 9;
         when "1100111000101" => index <= 8;
         when "1100111000110" => index <= 8;
         when "1100111000111" => index <= 7;
         when "1100111001000" => index <= 9;
         when "1100111001001" => index <= 8;
         when "1100111001010" => index <= 8;
         when "1100111001011" => index <= 7;
         when "1100111001100" => index <= 8;
         when "1100111001101" => index <= 7;
         when "1100111001110" => index <= 7;
         when "1100111001111" => index <= 7;
         when "1100111010000" => index <= 9;
         when "1100111010001" => index <= 8;
         when "1100111010010" => index <= 8;
         when "1100111010011" => index <= 7;
         when "1100111010100" => index <= 8;
         when "1100111010101" => index <= 7;
         when "1100111010110" => index <= 7;
         when "1100111010111" => index <= 7;
         when "1100111011000" => index <= 8;
         when "1100111011001" => index <= 7;
         when "1100111011010" => index <= 8;
         when "1100111011011" => index <= 7;
         when "1100111011100" => index <= 8;
         when "1100111011101" => index <= 7;
         when "1100111011110" => index <= 7;
         when "1100111011111" => index <= 6;
         when "1100111100000" => index <= 9;
         when "1100111100001" => index <= 8;
         when "1100111100010" => index <= 8;
         when "1100111100011" => index <= 7;
         when "1100111100100" => index <= 8;
         when "1100111100101" => index <= 7;
         when "1100111100110" => index <= 8;
         when "1100111100111" => index <= 7;
         when "1100111101000" => index <= 8;
         when "1100111101001" => index <= 8;
         when "1100111101010" => index <= 8;
         when "1100111101011" => index <= 7;
         when "1100111101100" => index <= 8;
         when "1100111101101" => index <= 7;
         when "1100111101110" => index <= 7;
         when "1100111101111" => index <= 6;
         when "1100111110000" => index <= 9;
         when "1100111110001" => index <= 8;
         when "1100111110010" => index <= 8;
         when "1100111110011" => index <= 7;
         when "1100111110100" => index <= 8;
         when "1100111110101" => index <= 7;
         when "1100111110110" => index <= 7;
         when "1100111110111" => index <= 7;
         when "1100111111000" => index <= 8;
         when "1100111111001" => index <= 7;
         when "1100111111010" => index <= 7;
         when "1100111111011" => index <= 7;
         when "1100111111100" => index <= 7;
         when "1100111111101" => index <= 7;
         when "1100111111110" => index <= 7;
         when "1100111111111" => index <= 6;
         when "1101000000000" => index <= 12;
         when "1101000000001" => index <= 9;
         when "1101000000010" => index <= 9;
         when "1101000000011" => index <= 8;
         when "1101000000100" => index <= 10;
         when "1101000000101" => index <= 8;
         when "1101000000110" => index <= 8;
         when "1101000000111" => index <= 7;
         when "1101000001000" => index <= 10;
         when "1101000001001" => index <= 8;
         when "1101000001010" => index <= 8;
         when "1101000001011" => index <= 7;
         when "1101000001100" => index <= 8;
         when "1101000001101" => index <= 7;
         when "1101000001110" => index <= 7;
         when "1101000001111" => index <= 6;
         when "1101000010000" => index <= 10;
         when "1101000010001" => index <= 8;
         when "1101000010010" => index <= 8;
         when "1101000010011" => index <= 7;
         when "1101000010100" => index <= 9;
         when "1101000010101" => index <= 7;
         when "1101000010110" => index <= 8;
         when "1101000010111" => index <= 7;
         when "1101000011000" => index <= 9;
         when "1101000011001" => index <= 8;
         when "1101000011010" => index <= 8;
         when "1101000011011" => index <= 7;
         when "1101000011100" => index <= 8;
         when "1101000011101" => index <= 7;
         when "1101000011110" => index <= 7;
         when "1101000011111" => index <= 6;
         when "1101000100000" => index <= 10;
         when "1101000100001" => index <= 8;
         when "1101000100010" => index <= 9;
         when "1101000100011" => index <= 7;
         when "1101000100100" => index <= 9;
         when "1101000100101" => index <= 8;
         when "1101000100110" => index <= 8;
         when "1101000100111" => index <= 7;
         when "1101000101000" => index <= 9;
         when "1101000101001" => index <= 8;
         when "1101000101010" => index <= 8;
         when "1101000101011" => index <= 7;
         when "1101000101100" => index <= 8;
         when "1101000101101" => index <= 7;
         when "1101000101110" => index <= 7;
         when "1101000101111" => index <= 6;
         when "1101000110000" => index <= 9;
         when "1101000110001" => index <= 8;
         when "1101000110010" => index <= 8;
         when "1101000110011" => index <= 7;
         when "1101000110100" => index <= 8;
         when "1101000110101" => index <= 7;
         when "1101000110110" => index <= 7;
         when "1101000110111" => index <= 6;
         when "1101000111000" => index <= 8;
         when "1101000111001" => index <= 7;
         when "1101000111010" => index <= 7;
         when "1101000111011" => index <= 7;
         when "1101000111100" => index <= 8;
         when "1101000111101" => index <= 7;
         when "1101000111110" => index <= 7;
         when "1101000111111" => index <= 6;
         when "1101001000000" => index <= 10;
         when "1101001000001" => index <= 9;
         when "1101001000010" => index <= 9;
         when "1101001000011" => index <= 8;
         when "1101001000100" => index <= 9;
         when "1101001000101" => index <= 8;
         when "1101001000110" => index <= 8;
         when "1101001000111" => index <= 7;
         when "1101001001000" => index <= 9;
         when "1101001001001" => index <= 8;
         when "1101001001010" => index <= 8;
         when "1101001001011" => index <= 7;
         when "1101001001100" => index <= 8;
         when "1101001001101" => index <= 7;
         when "1101001001110" => index <= 7;
         when "1101001001111" => index <= 6;
         when "1101001010000" => index <= 9;
         when "1101001010001" => index <= 8;
         when "1101001010010" => index <= 8;
         when "1101001010011" => index <= 7;
         when "1101001010100" => index <= 8;
         when "1101001010101" => index <= 7;
         when "1101001010110" => index <= 7;
         when "1101001010111" => index <= 7;
         when "1101001011000" => index <= 8;
         when "1101001011001" => index <= 7;
         when "1101001011010" => index <= 8;
         when "1101001011011" => index <= 7;
         when "1101001011100" => index <= 8;
         when "1101001011101" => index <= 7;
         when "1101001011110" => index <= 7;
         when "1101001011111" => index <= 6;
         when "1101001100000" => index <= 10;
         when "1101001100001" => index <= 8;
         when "1101001100010" => index <= 8;
         when "1101001100011" => index <= 7;
         when "1101001100100" => index <= 8;
         when "1101001100101" => index <= 7;
         when "1101001100110" => index <= 8;
         when "1101001100111" => index <= 7;
         when "1101001101000" => index <= 9;
         when "1101001101001" => index <= 8;
         when "1101001101010" => index <= 8;
         when "1101001101011" => index <= 7;
         when "1101001101100" => index <= 8;
         when "1101001101101" => index <= 7;
         when "1101001101110" => index <= 7;
         when "1101001101111" => index <= 6;
         when "1101001110000" => index <= 9;
         when "1101001110001" => index <= 8;
         when "1101001110010" => index <= 8;
         when "1101001110011" => index <= 7;
         when "1101001110100" => index <= 8;
         when "1101001110101" => index <= 7;
         when "1101001110110" => index <= 7;
         when "1101001110111" => index <= 7;
         when "1101001111000" => index <= 8;
         when "1101001111001" => index <= 7;
         when "1101001111010" => index <= 7;
         when "1101001111011" => index <= 7;
         when "1101001111100" => index <= 8;
         when "1101001111101" => index <= 7;
         when "1101001111110" => index <= 7;
         when "1101001111111" => index <= 6;
         when "1101010000000" => index <= 11;
         when "1101010000001" => index <= 9;
         when "1101010000010" => index <= 9;
         when "1101010000011" => index <= 8;
         when "1101010000100" => index <= 9;
         when "1101010000101" => index <= 8;
         when "1101010000110" => index <= 8;
         when "1101010000111" => index <= 7;
         when "1101010001000" => index <= 9;
         when "1101010001001" => index <= 8;
         when "1101010001010" => index <= 8;
         when "1101010001011" => index <= 7;
         when "1101010001100" => index <= 8;
         when "1101010001101" => index <= 7;
         when "1101010001110" => index <= 7;
         when "1101010001111" => index <= 7;
         when "1101010010000" => index <= 10;
         when "1101010010001" => index <= 8;
         when "1101010010010" => index <= 8;
         when "1101010010011" => index <= 7;
         when "1101010010100" => index <= 8;
         when "1101010010101" => index <= 7;
         when "1101010010110" => index <= 8;
         when "1101010010111" => index <= 7;
         when "1101010011000" => index <= 9;
         when "1101010011001" => index <= 8;
         when "1101010011010" => index <= 8;
         when "1101010011011" => index <= 7;
         when "1101010011100" => index <= 8;
         when "1101010011101" => index <= 7;
         when "1101010011110" => index <= 7;
         when "1101010011111" => index <= 6;
         when "1101010100000" => index <= 10;
         when "1101010100001" => index <= 8;
         when "1101010100010" => index <= 8;
         when "1101010100011" => index <= 7;
         when "1101010100100" => index <= 9;
         when "1101010100101" => index <= 8;
         when "1101010100110" => index <= 8;
         when "1101010100111" => index <= 7;
         when "1101010101000" => index <= 9;
         when "1101010101001" => index <= 8;
         when "1101010101010" => index <= 8;
         when "1101010101011" => index <= 7;
         when "1101010101100" => index <= 8;
         when "1101010101101" => index <= 7;
         when "1101010101110" => index <= 7;
         when "1101010101111" => index <= 7;
         when "1101010110000" => index <= 9;
         when "1101010110001" => index <= 8;
         when "1101010110010" => index <= 8;
         when "1101010110011" => index <= 7;
         when "1101010110100" => index <= 8;
         when "1101010110101" => index <= 7;
         when "1101010110110" => index <= 7;
         when "1101010110111" => index <= 7;
         when "1101010111000" => index <= 8;
         when "1101010111001" => index <= 7;
         when "1101010111010" => index <= 8;
         when "1101010111011" => index <= 7;
         when "1101010111100" => index <= 8;
         when "1101010111101" => index <= 7;
         when "1101010111110" => index <= 7;
         when "1101010111111" => index <= 6;
         when "1101011000000" => index <= 10;
         when "1101011000001" => index <= 8;
         when "1101011000010" => index <= 9;
         when "1101011000011" => index <= 8;
         when "1101011000100" => index <= 9;
         when "1101011000101" => index <= 8;
         when "1101011000110" => index <= 8;
         when "1101011000111" => index <= 7;
         when "1101011001000" => index <= 9;
         when "1101011001001" => index <= 8;
         when "1101011001010" => index <= 8;
         when "1101011001011" => index <= 7;
         when "1101011001100" => index <= 8;
         when "1101011001101" => index <= 7;
         when "1101011001110" => index <= 7;
         when "1101011001111" => index <= 7;
         when "1101011010000" => index <= 9;
         when "1101011010001" => index <= 8;
         when "1101011010010" => index <= 8;
         when "1101011010011" => index <= 7;
         when "1101011010100" => index <= 8;
         when "1101011010101" => index <= 7;
         when "1101011010110" => index <= 8;
         when "1101011010111" => index <= 7;
         when "1101011011000" => index <= 8;
         when "1101011011001" => index <= 8;
         when "1101011011010" => index <= 8;
         when "1101011011011" => index <= 7;
         when "1101011011100" => index <= 8;
         when "1101011011101" => index <= 7;
         when "1101011011110" => index <= 7;
         when "1101011011111" => index <= 6;
         when "1101011100000" => index <= 9;
         when "1101011100001" => index <= 8;
         when "1101011100010" => index <= 8;
         when "1101011100011" => index <= 7;
         when "1101011100100" => index <= 8;
         when "1101011100101" => index <= 8;
         when "1101011100110" => index <= 8;
         when "1101011100111" => index <= 7;
         when "1101011101000" => index <= 9;
         when "1101011101001" => index <= 8;
         when "1101011101010" => index <= 8;
         when "1101011101011" => index <= 7;
         when "1101011101100" => index <= 8;
         when "1101011101101" => index <= 7;
         when "1101011101110" => index <= 7;
         when "1101011101111" => index <= 7;
         when "1101011110000" => index <= 9;
         when "1101011110001" => index <= 8;
         when "1101011110010" => index <= 8;
         when "1101011110011" => index <= 7;
         when "1101011110100" => index <= 8;
         when "1101011110101" => index <= 7;
         when "1101011110110" => index <= 7;
         when "1101011110111" => index <= 7;
         when "1101011111000" => index <= 8;
         when "1101011111001" => index <= 7;
         when "1101011111010" => index <= 7;
         when "1101011111011" => index <= 7;
         when "1101011111100" => index <= 8;
         when "1101011111101" => index <= 7;
         when "1101011111110" => index <= 7;
         when "1101011111111" => index <= 6;
         when "1101100000000" => index <= 11;
         when "1101100000001" => index <= 9;
         when "1101100000010" => index <= 9;
         when "1101100000011" => index <= 8;
         when "1101100000100" => index <= 9;
         when "1101100000101" => index <= 8;
         when "1101100000110" => index <= 8;
         when "1101100000111" => index <= 7;
         when "1101100001000" => index <= 10;
         when "1101100001001" => index <= 8;
         when "1101100001010" => index <= 8;
         when "1101100001011" => index <= 7;
         when "1101100001100" => index <= 8;
         when "1101100001101" => index <= 7;
         when "1101100001110" => index <= 8;
         when "1101100001111" => index <= 7;
         when "1101100010000" => index <= 10;
         when "1101100010001" => index <= 8;
         when "1101100010010" => index <= 8;
         when "1101100010011" => index <= 7;
         when "1101100010100" => index <= 9;
         when "1101100010101" => index <= 8;
         when "1101100010110" => index <= 8;
         when "1101100010111" => index <= 7;
         when "1101100011000" => index <= 9;
         when "1101100011001" => index <= 8;
         when "1101100011010" => index <= 8;
         when "1101100011011" => index <= 7;
         when "1101100011100" => index <= 8;
         when "1101100011101" => index <= 7;
         when "1101100011110" => index <= 7;
         when "1101100011111" => index <= 7;
         when "1101100100000" => index <= 10;
         when "1101100100001" => index <= 8;
         when "1101100100010" => index <= 9;
         when "1101100100011" => index <= 8;
         when "1101100100100" => index <= 9;
         when "1101100100101" => index <= 8;
         when "1101100100110" => index <= 8;
         when "1101100100111" => index <= 7;
         when "1101100101000" => index <= 9;
         when "1101100101001" => index <= 8;
         when "1101100101010" => index <= 8;
         when "1101100101011" => index <= 7;
         when "1101100101100" => index <= 8;
         when "1101100101101" => index <= 7;
         when "1101100101110" => index <= 7;
         when "1101100101111" => index <= 7;
         when "1101100110000" => index <= 9;
         when "1101100110001" => index <= 8;
         when "1101100110010" => index <= 8;
         when "1101100110011" => index <= 7;
         when "1101100110100" => index <= 8;
         when "1101100110101" => index <= 7;
         when "1101100110110" => index <= 8;
         when "1101100110111" => index <= 7;
         when "1101100111000" => index <= 8;
         when "1101100111001" => index <= 8;
         when "1101100111010" => index <= 8;
         when "1101100111011" => index <= 7;
         when "1101100111100" => index <= 8;
         when "1101100111101" => index <= 7;
         when "1101100111110" => index <= 7;
         when "1101100111111" => index <= 6;
         when "1101101000000" => index <= 10;
         when "1101101000001" => index <= 9;
         when "1101101000010" => index <= 9;
         when "1101101000011" => index <= 8;
         when "1101101000100" => index <= 9;
         when "1101101000101" => index <= 8;
         when "1101101000110" => index <= 8;
         when "1101101000111" => index <= 7;
         when "1101101001000" => index <= 9;
         when "1101101001001" => index <= 8;
         when "1101101001010" => index <= 8;
         when "1101101001011" => index <= 7;
         when "1101101001100" => index <= 8;
         when "1101101001101" => index <= 7;
         when "1101101001110" => index <= 8;
         when "1101101001111" => index <= 7;
         when "1101101010000" => index <= 9;
         when "1101101010001" => index <= 8;
         when "1101101010010" => index <= 8;
         when "1101101010011" => index <= 7;
         when "1101101010100" => index <= 8;
         when "1101101010101" => index <= 8;
         when "1101101010110" => index <= 8;
         when "1101101010111" => index <= 7;
         when "1101101011000" => index <= 9;
         when "1101101011001" => index <= 8;
         when "1101101011010" => index <= 8;
         when "1101101011011" => index <= 7;
         when "1101101011100" => index <= 8;
         when "1101101011101" => index <= 7;
         when "1101101011110" => index <= 7;
         when "1101101011111" => index <= 7;
         when "1101101100000" => index <= 10;
         when "1101101100001" => index <= 8;
         when "1101101100010" => index <= 8;
         when "1101101100011" => index <= 8;
         when "1101101100100" => index <= 9;
         when "1101101100101" => index <= 8;
         when "1101101100110" => index <= 8;
         when "1101101100111" => index <= 7;
         when "1101101101000" => index <= 9;
         when "1101101101001" => index <= 8;
         when "1101101101010" => index <= 8;
         when "1101101101011" => index <= 7;
         when "1101101101100" => index <= 8;
         when "1101101101101" => index <= 7;
         when "1101101101110" => index <= 7;
         when "1101101101111" => index <= 7;
         when "1101101110000" => index <= 9;
         when "1101101110001" => index <= 8;
         when "1101101110010" => index <= 8;
         when "1101101110011" => index <= 7;
         when "1101101110100" => index <= 8;
         when "1101101110101" => index <= 7;
         when "1101101110110" => index <= 7;
         when "1101101110111" => index <= 7;
         when "1101101111000" => index <= 8;
         when "1101101111001" => index <= 7;
         when "1101101111010" => index <= 8;
         when "1101101111011" => index <= 7;
         when "1101101111100" => index <= 8;
         when "1101101111101" => index <= 7;
         when "1101101111110" => index <= 7;
         when "1101101111111" => index <= 7;
         when "1101110000000" => index <= 10;
         when "1101110000001" => index <= 9;
         when "1101110000010" => index <= 9;
         when "1101110000011" => index <= 8;
         when "1101110000100" => index <= 9;
         when "1101110000101" => index <= 8;
         when "1101110000110" => index <= 8;
         when "1101110000111" => index <= 7;
         when "1101110001000" => index <= 9;
         when "1101110001001" => index <= 8;
         when "1101110001010" => index <= 8;
         when "1101110001011" => index <= 7;
         when "1101110001100" => index <= 8;
         when "1101110001101" => index <= 8;
         when "1101110001110" => index <= 8;
         when "1101110001111" => index <= 7;
         when "1101110010000" => index <= 10;
         when "1101110010001" => index <= 8;
         when "1101110010010" => index <= 8;
         when "1101110010011" => index <= 8;
         when "1101110010100" => index <= 9;
         when "1101110010101" => index <= 8;
         when "1101110010110" => index <= 8;
         when "1101110010111" => index <= 7;
         when "1101110011000" => index <= 9;
         when "1101110011001" => index <= 8;
         when "1101110011010" => index <= 8;
         when "1101110011011" => index <= 7;
         when "1101110011100" => index <= 8;
         when "1101110011101" => index <= 7;
         when "1101110011110" => index <= 7;
         when "1101110011111" => index <= 7;
         when "1101110100000" => index <= 10;
         when "1101110100001" => index <= 8;
         when "1101110100010" => index <= 9;
         when "1101110100011" => index <= 8;
         when "1101110100100" => index <= 9;
         when "1101110100101" => index <= 8;
         when "1101110100110" => index <= 8;
         when "1101110100111" => index <= 7;
         when "1101110101000" => index <= 9;
         when "1101110101001" => index <= 8;
         when "1101110101010" => index <= 8;
         when "1101110101011" => index <= 7;
         when "1101110101100" => index <= 8;
         when "1101110101101" => index <= 7;
         when "1101110101110" => index <= 7;
         when "1101110101111" => index <= 7;
         when "1101110110000" => index <= 9;
         when "1101110110001" => index <= 8;
         when "1101110110010" => index <= 8;
         when "1101110110011" => index <= 7;
         when "1101110110100" => index <= 8;
         when "1101110110101" => index <= 7;
         when "1101110110110" => index <= 8;
         when "1101110110111" => index <= 7;
         when "1101110111000" => index <= 8;
         when "1101110111001" => index <= 8;
         when "1101110111010" => index <= 8;
         when "1101110111011" => index <= 7;
         when "1101110111100" => index <= 8;
         when "1101110111101" => index <= 7;
         when "1101110111110" => index <= 7;
         when "1101110111111" => index <= 7;
         when "1101111000000" => index <= 10;
         when "1101111000001" => index <= 9;
         when "1101111000010" => index <= 9;
         when "1101111000011" => index <= 8;
         when "1101111000100" => index <= 9;
         when "1101111000101" => index <= 8;
         when "1101111000110" => index <= 8;
         when "1101111000111" => index <= 7;
         when "1101111001000" => index <= 9;
         when "1101111001001" => index <= 8;
         when "1101111001010" => index <= 8;
         when "1101111001011" => index <= 7;
         when "1101111001100" => index <= 8;
         when "1101111001101" => index <= 7;
         when "1101111001110" => index <= 8;
         when "1101111001111" => index <= 7;
         when "1101111010000" => index <= 9;
         when "1101111010001" => index <= 8;
         when "1101111010010" => index <= 8;
         when "1101111010011" => index <= 7;
         when "1101111010100" => index <= 8;
         when "1101111010101" => index <= 8;
         when "1101111010110" => index <= 8;
         when "1101111010111" => index <= 7;
         when "1101111011000" => index <= 8;
         when "1101111011001" => index <= 8;
         when "1101111011010" => index <= 8;
         when "1101111011011" => index <= 7;
         when "1101111011100" => index <= 8;
         when "1101111011101" => index <= 7;
         when "1101111011110" => index <= 7;
         when "1101111011111" => index <= 7;
         when "1101111100000" => index <= 9;
         when "1101111100001" => index <= 8;
         when "1101111100010" => index <= 8;
         when "1101111100011" => index <= 8;
         when "1101111100100" => index <= 8;
         when "1101111100101" => index <= 8;
         when "1101111100110" => index <= 8;
         when "1101111100111" => index <= 7;
         when "1101111101000" => index <= 9;
         when "1101111101001" => index <= 8;
         when "1101111101010" => index <= 8;
         when "1101111101011" => index <= 7;
         when "1101111101100" => index <= 8;
         when "1101111101101" => index <= 7;
         when "1101111101110" => index <= 7;
         when "1101111101111" => index <= 7;
         when "1101111110000" => index <= 9;
         when "1101111110001" => index <= 8;
         when "1101111110010" => index <= 8;
         when "1101111110011" => index <= 7;
         when "1101111110100" => index <= 8;
         when "1101111110101" => index <= 7;
         when "1101111110110" => index <= 8;
         when "1101111110111" => index <= 7;
         when "1101111111000" => index <= 8;
         when "1101111111001" => index <= 8;
         when "1101111111010" => index <= 8;
         when "1101111111011" => index <= 7;
         when "1101111111100" => index <= 8;
         when "1101111111101" => index <= 7;
         when "1101111111110" => index <= 7;
         when "1101111111111" => index <= 7;
         when "1110000000000" => index <= 12;
         when "1110000000001" => index <= 9;
         when "1110000000010" => index <= 10;
         when "1110000000011" => index <= 8;
         when "1110000000100" => index <= 10;
         when "1110000000101" => index <= 8;
         when "1110000000110" => index <= 8;
         when "1110000000111" => index <= 7;
         when "1110000001000" => index <= 10;
         when "1110000001001" => index <= 8;
         when "1110000001010" => index <= 8;
         when "1110000001011" => index <= 7;
         when "1110000001100" => index <= 9;
         when "1110000001101" => index <= 7;
         when "1110000001110" => index <= 8;
         when "1110000001111" => index <= 7;
         when "1110000010000" => index <= 10;
         when "1110000010001" => index <= 8;
         when "1110000010010" => index <= 9;
         when "1110000010011" => index <= 7;
         when "1110000010100" => index <= 9;
         when "1110000010101" => index <= 8;
         when "1110000010110" => index <= 8;
         when "1110000010111" => index <= 7;
         when "1110000011000" => index <= 9;
         when "1110000011001" => index <= 8;
         when "1110000011010" => index <= 8;
         when "1110000011011" => index <= 7;
         when "1110000011100" => index <= 8;
         when "1110000011101" => index <= 7;
         when "1110000011110" => index <= 7;
         when "1110000011111" => index <= 6;
         when "1110000100000" => index <= 10;
         when "1110000100001" => index <= 9;
         when "1110000100010" => index <= 9;
         when "1110000100011" => index <= 8;
         when "1110000100100" => index <= 9;
         when "1110000100101" => index <= 8;
         when "1110000100110" => index <= 8;
         when "1110000100111" => index <= 7;
         when "1110000101000" => index <= 9;
         when "1110000101001" => index <= 8;
         when "1110000101010" => index <= 8;
         when "1110000101011" => index <= 7;
         when "1110000101100" => index <= 8;
         when "1110000101101" => index <= 7;
         when "1110000101110" => index <= 7;
         when "1110000101111" => index <= 6;
         when "1110000110000" => index <= 9;
         when "1110000110001" => index <= 8;
         when "1110000110010" => index <= 8;
         when "1110000110011" => index <= 7;
         when "1110000110100" => index <= 8;
         when "1110000110101" => index <= 7;
         when "1110000110110" => index <= 7;
         when "1110000110111" => index <= 7;
         when "1110000111000" => index <= 8;
         when "1110000111001" => index <= 7;
         when "1110000111010" => index <= 8;
         when "1110000111011" => index <= 7;
         when "1110000111100" => index <= 8;
         when "1110000111101" => index <= 7;
         when "1110000111110" => index <= 7;
         when "1110000111111" => index <= 6;
         when "1110001000000" => index <= 11;
         when "1110001000001" => index <= 9;
         when "1110001000010" => index <= 9;
         when "1110001000011" => index <= 8;
         when "1110001000100" => index <= 9;
         when "1110001000101" => index <= 8;
         when "1110001000110" => index <= 8;
         when "1110001000111" => index <= 7;
         when "1110001001000" => index <= 9;
         when "1110001001001" => index <= 8;
         when "1110001001010" => index <= 8;
         when "1110001001011" => index <= 7;
         when "1110001001100" => index <= 8;
         when "1110001001101" => index <= 7;
         when "1110001001110" => index <= 7;
         when "1110001001111" => index <= 7;
         when "1110001010000" => index <= 10;
         when "1110001010001" => index <= 8;
         when "1110001010010" => index <= 8;
         when "1110001010011" => index <= 7;
         when "1110001010100" => index <= 8;
         when "1110001010101" => index <= 7;
         when "1110001010110" => index <= 8;
         when "1110001010111" => index <= 7;
         when "1110001011000" => index <= 9;
         when "1110001011001" => index <= 8;
         when "1110001011010" => index <= 8;
         when "1110001011011" => index <= 7;
         when "1110001011100" => index <= 8;
         when "1110001011101" => index <= 7;
         when "1110001011110" => index <= 7;
         when "1110001011111" => index <= 6;
         when "1110001100000" => index <= 10;
         when "1110001100001" => index <= 8;
         when "1110001100010" => index <= 8;
         when "1110001100011" => index <= 7;
         when "1110001100100" => index <= 9;
         when "1110001100101" => index <= 8;
         when "1110001100110" => index <= 8;
         when "1110001100111" => index <= 7;
         when "1110001101000" => index <= 9;
         when "1110001101001" => index <= 8;
         when "1110001101010" => index <= 8;
         when "1110001101011" => index <= 7;
         when "1110001101100" => index <= 8;
         when "1110001101101" => index <= 7;
         when "1110001101110" => index <= 7;
         when "1110001101111" => index <= 7;
         when "1110001110000" => index <= 9;
         when "1110001110001" => index <= 8;
         when "1110001110010" => index <= 8;
         when "1110001110011" => index <= 7;
         when "1110001110100" => index <= 8;
         when "1110001110101" => index <= 7;
         when "1110001110110" => index <= 7;
         when "1110001110111" => index <= 7;
         when "1110001111000" => index <= 8;
         when "1110001111001" => index <= 7;
         when "1110001111010" => index <= 8;
         when "1110001111011" => index <= 7;
         when "1110001111100" => index <= 8;
         when "1110001111101" => index <= 7;
         when "1110001111110" => index <= 7;
         when "1110001111111" => index <= 6;
         when "1110010000000" => index <= 11;
         when "1110010000001" => index <= 9;
         when "1110010000010" => index <= 9;
         when "1110010000011" => index <= 8;
         when "1110010000100" => index <= 9;
         when "1110010000101" => index <= 8;
         when "1110010000110" => index <= 8;
         when "1110010000111" => index <= 7;
         when "1110010001000" => index <= 10;
         when "1110010001001" => index <= 8;
         when "1110010001010" => index <= 8;
         when "1110010001011" => index <= 7;
         when "1110010001100" => index <= 8;
         when "1110010001101" => index <= 7;
         when "1110010001110" => index <= 8;
         when "1110010001111" => index <= 7;
         when "1110010010000" => index <= 10;
         when "1110010010001" => index <= 8;
         when "1110010010010" => index <= 8;
         when "1110010010011" => index <= 7;
         when "1110010010100" => index <= 9;
         when "1110010010101" => index <= 8;
         when "1110010010110" => index <= 8;
         when "1110010010111" => index <= 7;
         when "1110010011000" => index <= 9;
         when "1110010011001" => index <= 8;
         when "1110010011010" => index <= 8;
         when "1110010011011" => index <= 7;
         when "1110010011100" => index <= 8;
         when "1110010011101" => index <= 7;
         when "1110010011110" => index <= 7;
         when "1110010011111" => index <= 7;
         when "1110010100000" => index <= 10;
         when "1110010100001" => index <= 8;
         when "1110010100010" => index <= 9;
         when "1110010100011" => index <= 8;
         when "1110010100100" => index <= 9;
         when "1110010100101" => index <= 8;
         when "1110010100110" => index <= 8;
         when "1110010100111" => index <= 7;
         when "1110010101000" => index <= 9;
         when "1110010101001" => index <= 8;
         when "1110010101010" => index <= 8;
         when "1110010101011" => index <= 7;
         when "1110010101100" => index <= 8;
         when "1110010101101" => index <= 7;
         when "1110010101110" => index <= 7;
         when "1110010101111" => index <= 7;
         when "1110010110000" => index <= 9;
         when "1110010110001" => index <= 8;
         when "1110010110010" => index <= 8;
         when "1110010110011" => index <= 7;
         when "1110010110100" => index <= 8;
         when "1110010110101" => index <= 7;
         when "1110010110110" => index <= 8;
         when "1110010110111" => index <= 7;
         when "1110010111000" => index <= 8;
         when "1110010111001" => index <= 8;
         when "1110010111010" => index <= 8;
         when "1110010111011" => index <= 7;
         when "1110010111100" => index <= 8;
         when "1110010111101" => index <= 7;
         when "1110010111110" => index <= 7;
         when "1110010111111" => index <= 6;
         when "1110011000000" => index <= 10;
         when "1110011000001" => index <= 9;
         when "1110011000010" => index <= 9;
         when "1110011000011" => index <= 8;
         when "1110011000100" => index <= 9;
         when "1110011000101" => index <= 8;
         when "1110011000110" => index <= 8;
         when "1110011000111" => index <= 7;
         when "1110011001000" => index <= 9;
         when "1110011001001" => index <= 8;
         when "1110011001010" => index <= 8;
         when "1110011001011" => index <= 7;
         when "1110011001100" => index <= 8;
         when "1110011001101" => index <= 7;
         when "1110011001110" => index <= 8;
         when "1110011001111" => index <= 7;
         when "1110011010000" => index <= 9;
         when "1110011010001" => index <= 8;
         when "1110011010010" => index <= 8;
         when "1110011010011" => index <= 7;
         when "1110011010100" => index <= 8;
         when "1110011010101" => index <= 8;
         when "1110011010110" => index <= 8;
         when "1110011010111" => index <= 7;
         when "1110011011000" => index <= 9;
         when "1110011011001" => index <= 8;
         when "1110011011010" => index <= 8;
         when "1110011011011" => index <= 7;
         when "1110011011100" => index <= 8;
         when "1110011011101" => index <= 7;
         when "1110011011110" => index <= 7;
         when "1110011011111" => index <= 7;
         when "1110011100000" => index <= 10;
         when "1110011100001" => index <= 8;
         when "1110011100010" => index <= 8;
         when "1110011100011" => index <= 8;
         when "1110011100100" => index <= 9;
         when "1110011100101" => index <= 8;
         when "1110011100110" => index <= 8;
         when "1110011100111" => index <= 7;
         when "1110011101000" => index <= 9;
         when "1110011101001" => index <= 8;
         when "1110011101010" => index <= 8;
         when "1110011101011" => index <= 7;
         when "1110011101100" => index <= 8;
         when "1110011101101" => index <= 7;
         when "1110011101110" => index <= 7;
         when "1110011101111" => index <= 7;
         when "1110011110000" => index <= 9;
         when "1110011110001" => index <= 8;
         when "1110011110010" => index <= 8;
         when "1110011110011" => index <= 7;
         when "1110011110100" => index <= 8;
         when "1110011110101" => index <= 7;
         when "1110011110110" => index <= 7;
         when "1110011110111" => index <= 7;
         when "1110011111000" => index <= 8;
         when "1110011111001" => index <= 7;
         when "1110011111010" => index <= 8;
         when "1110011111011" => index <= 7;
         when "1110011111100" => index <= 8;
         when "1110011111101" => index <= 7;
         when "1110011111110" => index <= 7;
         when "1110011111111" => index <= 7;
         when "1110100000000" => index <= 11;
         when "1110100000001" => index <= 9;
         when "1110100000010" => index <= 9;
         when "1110100000011" => index <= 8;
         when "1110100000100" => index <= 10;
         when "1110100000101" => index <= 8;
         when "1110100000110" => index <= 8;
         when "1110100000111" => index <= 7;
         when "1110100001000" => index <= 10;
         when "1110100001001" => index <= 8;
         when "1110100001010" => index <= 8;
         when "1110100001011" => index <= 7;
         when "1110100001100" => index <= 9;
         when "1110100001101" => index <= 8;
         when "1110100001110" => index <= 8;
         when "1110100001111" => index <= 7;
         when "1110100010000" => index <= 10;
         when "1110100010001" => index <= 8;
         when "1110100010010" => index <= 9;
         when "1110100010011" => index <= 8;
         when "1110100010100" => index <= 9;
         when "1110100010101" => index <= 8;
         when "1110100010110" => index <= 8;
         when "1110100010111" => index <= 7;
         when "1110100011000" => index <= 9;
         when "1110100011001" => index <= 8;
         when "1110100011010" => index <= 8;
         when "1110100011011" => index <= 7;
         when "1110100011100" => index <= 8;
         when "1110100011101" => index <= 7;
         when "1110100011110" => index <= 7;
         when "1110100011111" => index <= 7;
         when "1110100100000" => index <= 10;
         when "1110100100001" => index <= 9;
         when "1110100100010" => index <= 9;
         when "1110100100011" => index <= 8;
         when "1110100100100" => index <= 9;
         when "1110100100101" => index <= 8;
         when "1110100100110" => index <= 8;
         when "1110100100111" => index <= 7;
         when "1110100101000" => index <= 9;
         when "1110100101001" => index <= 8;
         when "1110100101010" => index <= 8;
         when "1110100101011" => index <= 7;
         when "1110100101100" => index <= 8;
         when "1110100101101" => index <= 7;
         when "1110100101110" => index <= 8;
         when "1110100101111" => index <= 7;
         when "1110100110000" => index <= 9;
         when "1110100110001" => index <= 8;
         when "1110100110010" => index <= 8;
         when "1110100110011" => index <= 7;
         when "1110100110100" => index <= 8;
         when "1110100110101" => index <= 8;
         when "1110100110110" => index <= 8;
         when "1110100110111" => index <= 7;
         when "1110100111000" => index <= 9;
         when "1110100111001" => index <= 8;
         when "1110100111010" => index <= 8;
         when "1110100111011" => index <= 7;
         when "1110100111100" => index <= 8;
         when "1110100111101" => index <= 7;
         when "1110100111110" => index <= 7;
         when "1110100111111" => index <= 7;
         when "1110101000000" => index <= 10;
         when "1110101000001" => index <= 9;
         when "1110101000010" => index <= 9;
         when "1110101000011" => index <= 8;
         when "1110101000100" => index <= 9;
         when "1110101000101" => index <= 8;
         when "1110101000110" => index <= 8;
         when "1110101000111" => index <= 7;
         when "1110101001000" => index <= 9;
         when "1110101001001" => index <= 8;
         when "1110101001010" => index <= 8;
         when "1110101001011" => index <= 7;
         when "1110101001100" => index <= 8;
         when "1110101001101" => index <= 8;
         when "1110101001110" => index <= 8;
         when "1110101001111" => index <= 7;
         when "1110101010000" => index <= 10;
         when "1110101010001" => index <= 8;
         when "1110101010010" => index <= 8;
         when "1110101010011" => index <= 8;
         when "1110101010100" => index <= 9;
         when "1110101010101" => index <= 8;
         when "1110101010110" => index <= 8;
         when "1110101010111" => index <= 7;
         when "1110101011000" => index <= 9;
         when "1110101011001" => index <= 8;
         when "1110101011010" => index <= 8;
         when "1110101011011" => index <= 7;
         when "1110101011100" => index <= 8;
         when "1110101011101" => index <= 7;
         when "1110101011110" => index <= 7;
         when "1110101011111" => index <= 7;
         when "1110101100000" => index <= 10;
         when "1110101100001" => index <= 8;
         when "1110101100010" => index <= 9;
         when "1110101100011" => index <= 8;
         when "1110101100100" => index <= 9;
         when "1110101100101" => index <= 8;
         when "1110101100110" => index <= 8;
         when "1110101100111" => index <= 7;
         when "1110101101000" => index <= 9;
         when "1110101101001" => index <= 8;
         when "1110101101010" => index <= 8;
         when "1110101101011" => index <= 7;
         when "1110101101100" => index <= 8;
         when "1110101101101" => index <= 7;
         when "1110101101110" => index <= 7;
         when "1110101101111" => index <= 7;
         when "1110101110000" => index <= 9;
         when "1110101110001" => index <= 8;
         when "1110101110010" => index <= 8;
         when "1110101110011" => index <= 7;
         when "1110101110100" => index <= 8;
         when "1110101110101" => index <= 7;
         when "1110101110110" => index <= 8;
         when "1110101110111" => index <= 7;
         when "1110101111000" => index <= 8;
         when "1110101111001" => index <= 8;
         when "1110101111010" => index <= 8;
         when "1110101111011" => index <= 7;
         when "1110101111100" => index <= 8;
         when "1110101111101" => index <= 7;
         when "1110101111110" => index <= 7;
         when "1110101111111" => index <= 7;
         when "1110110000000" => index <= 11;
         when "1110110000001" => index <= 9;
         when "1110110000010" => index <= 9;
         when "1110110000011" => index <= 8;
         when "1110110000100" => index <= 9;
         when "1110110000101" => index <= 8;
         when "1110110000110" => index <= 8;
         when "1110110000111" => index <= 7;
         when "1110110001000" => index <= 10;
         when "1110110001001" => index <= 8;
         when "1110110001010" => index <= 8;
         when "1110110001011" => index <= 8;
         when "1110110001100" => index <= 9;
         when "1110110001101" => index <= 8;
         when "1110110001110" => index <= 8;
         when "1110110001111" => index <= 7;
         when "1110110010000" => index <= 10;
         when "1110110010001" => index <= 8;
         when "1110110010010" => index <= 9;
         when "1110110010011" => index <= 8;
         when "1110110010100" => index <= 9;
         when "1110110010101" => index <= 8;
         when "1110110010110" => index <= 8;
         when "1110110010111" => index <= 7;
         when "1110110011000" => index <= 9;
         when "1110110011001" => index <= 8;
         when "1110110011010" => index <= 8;
         when "1110110011011" => index <= 7;
         when "1110110011100" => index <= 8;
         when "1110110011101" => index <= 7;
         when "1110110011110" => index <= 7;
         when "1110110011111" => index <= 7;
         when "1110110100000" => index <= 10;
         when "1110110100001" => index <= 9;
         when "1110110100010" => index <= 9;
         when "1110110100011" => index <= 8;
         when "1110110100100" => index <= 9;
         when "1110110100101" => index <= 8;
         when "1110110100110" => index <= 8;
         when "1110110100111" => index <= 7;
         when "1110110101000" => index <= 9;
         when "1110110101001" => index <= 8;
         when "1110110101010" => index <= 8;
         when "1110110101011" => index <= 7;
         when "1110110101100" => index <= 8;
         when "1110110101101" => index <= 7;
         when "1110110101110" => index <= 8;
         when "1110110101111" => index <= 7;
         when "1110110110000" => index <= 9;
         when "1110110110001" => index <= 8;
         when "1110110110010" => index <= 8;
         when "1110110110011" => index <= 7;
         when "1110110110100" => index <= 8;
         when "1110110110101" => index <= 8;
         when "1110110110110" => index <= 8;
         when "1110110110111" => index <= 7;
         when "1110110111000" => index <= 8;
         when "1110110111001" => index <= 8;
         when "1110110111010" => index <= 8;
         when "1110110111011" => index <= 7;
         when "1110110111100" => index <= 8;
         when "1110110111101" => index <= 7;
         when "1110110111110" => index <= 7;
         when "1110110111111" => index <= 7;
         when "1110111000000" => index <= 10;
         when "1110111000001" => index <= 9;
         when "1110111000010" => index <= 9;
         when "1110111000011" => index <= 8;
         when "1110111000100" => index <= 9;
         when "1110111000101" => index <= 8;
         when "1110111000110" => index <= 8;
         when "1110111000111" => index <= 7;
         when "1110111001000" => index <= 9;
         when "1110111001001" => index <= 8;
         when "1110111001010" => index <= 8;
         when "1110111001011" => index <= 7;
         when "1110111001100" => index <= 8;
         when "1110111001101" => index <= 8;
         when "1110111001110" => index <= 8;
         when "1110111001111" => index <= 7;
         when "1110111010000" => index <= 9;
         when "1110111010001" => index <= 8;
         when "1110111010010" => index <= 8;
         when "1110111010011" => index <= 8;
         when "1110111010100" => index <= 8;
         when "1110111010101" => index <= 8;
         when "1110111010110" => index <= 8;
         when "1110111010111" => index <= 7;
         when "1110111011000" => index <= 9;
         when "1110111011001" => index <= 8;
         when "1110111011010" => index <= 8;
         when "1110111011011" => index <= 7;
         when "1110111011100" => index <= 8;
         when "1110111011101" => index <= 7;
         when "1110111011110" => index <= 7;
         when "1110111011111" => index <= 7;
         when "1110111100000" => index <= 9;
         when "1110111100001" => index <= 8;
         when "1110111100010" => index <= 8;
         when "1110111100011" => index <= 8;
         when "1110111100100" => index <= 9;
         when "1110111100101" => index <= 8;
         when "1110111100110" => index <= 8;
         when "1110111100111" => index <= 7;
         when "1110111101000" => index <= 9;
         when "1110111101001" => index <= 8;
         when "1110111101010" => index <= 8;
         when "1110111101011" => index <= 7;
         when "1110111101100" => index <= 8;
         when "1110111101101" => index <= 7;
         when "1110111101110" => index <= 8;
         when "1110111101111" => index <= 7;
         when "1110111110000" => index <= 9;
         when "1110111110001" => index <= 8;
         when "1110111110010" => index <= 8;
         when "1110111110011" => index <= 7;
         when "1110111110100" => index <= 8;
         when "1110111110101" => index <= 8;
         when "1110111110110" => index <= 8;
         when "1110111110111" => index <= 7;
         when "1110111111000" => index <= 8;
         when "1110111111001" => index <= 8;
         when "1110111111010" => index <= 8;
         when "1110111111011" => index <= 7;
         when "1110111111100" => index <= 8;
         when "1110111111101" => index <= 7;
         when "1110111111110" => index <= 7;
         when "1110111111111" => index <= 7;
         when "1111000000000" => index <= 12;
         when "1111000000001" => index <= 9;
         when "1111000000010" => index <= 10;
         when "1111000000011" => index <= 8;
         when "1111000000100" => index <= 10;
         when "1111000000101" => index <= 8;
         when "1111000000110" => index <= 8;
         when "1111000000111" => index <= 7;
         when "1111000001000" => index <= 10;
         when "1111000001001" => index <= 8;
         when "1111000001010" => index <= 9;
         when "1111000001011" => index <= 8;
         when "1111000001100" => index <= 9;
         when "1111000001101" => index <= 8;
         when "1111000001110" => index <= 8;
         when "1111000001111" => index <= 7;
         when "1111000010000" => index <= 10;
         when "1111000010001" => index <= 9;
         when "1111000010010" => index <= 9;
         when "1111000010011" => index <= 8;
         when "1111000010100" => index <= 9;
         when "1111000010101" => index <= 8;
         when "1111000010110" => index <= 8;
         when "1111000010111" => index <= 7;
         when "1111000011000" => index <= 9;
         when "1111000011001" => index <= 8;
         when "1111000011010" => index <= 8;
         when "1111000011011" => index <= 7;
         when "1111000011100" => index <= 8;
         when "1111000011101" => index <= 7;
         when "1111000011110" => index <= 8;
         when "1111000011111" => index <= 7;
         when "1111000100000" => index <= 10;
         when "1111000100001" => index <= 9;
         when "1111000100010" => index <= 9;
         when "1111000100011" => index <= 8;
         when "1111000100100" => index <= 9;
         when "1111000100101" => index <= 8;
         when "1111000100110" => index <= 8;
         when "1111000100111" => index <= 7;
         when "1111000101000" => index <= 9;
         when "1111000101001" => index <= 8;
         when "1111000101010" => index <= 8;
         when "1111000101011" => index <= 7;
         when "1111000101100" => index <= 8;
         when "1111000101101" => index <= 8;
         when "1111000101110" => index <= 8;
         when "1111000101111" => index <= 7;
         when "1111000110000" => index <= 10;
         when "1111000110001" => index <= 8;
         when "1111000110010" => index <= 8;
         when "1111000110011" => index <= 8;
         when "1111000110100" => index <= 9;
         when "1111000110101" => index <= 8;
         when "1111000110110" => index <= 8;
         when "1111000110111" => index <= 7;
         when "1111000111000" => index <= 9;
         when "1111000111001" => index <= 8;
         when "1111000111010" => index <= 8;
         when "1111000111011" => index <= 7;
         when "1111000111100" => index <= 8;
         when "1111000111101" => index <= 7;
         when "1111000111110" => index <= 7;
         when "1111000111111" => index <= 7;
         when "1111001000000" => index <= 11;
         when "1111001000001" => index <= 9;
         when "1111001000010" => index <= 9;
         when "1111001000011" => index <= 8;
         when "1111001000100" => index <= 9;
         when "1111001000101" => index <= 8;
         when "1111001000110" => index <= 8;
         when "1111001000111" => index <= 7;
         when "1111001001000" => index <= 10;
         when "1111001001001" => index <= 8;
         when "1111001001010" => index <= 8;
         when "1111001001011" => index <= 8;
         when "1111001001100" => index <= 9;
         when "1111001001101" => index <= 8;
         when "1111001001110" => index <= 8;
         when "1111001001111" => index <= 7;
         when "1111001010000" => index <= 10;
         when "1111001010001" => index <= 8;
         when "1111001010010" => index <= 9;
         when "1111001010011" => index <= 8;
         when "1111001010100" => index <= 9;
         when "1111001010101" => index <= 8;
         when "1111001010110" => index <= 8;
         when "1111001010111" => index <= 7;
         when "1111001011000" => index <= 9;
         when "1111001011001" => index <= 8;
         when "1111001011010" => index <= 8;
         when "1111001011011" => index <= 7;
         when "1111001011100" => index <= 8;
         when "1111001011101" => index <= 7;
         when "1111001011110" => index <= 7;
         when "1111001011111" => index <= 7;
         when "1111001100000" => index <= 10;
         when "1111001100001" => index <= 9;
         when "1111001100010" => index <= 9;
         when "1111001100011" => index <= 8;
         when "1111001100100" => index <= 9;
         when "1111001100101" => index <= 8;
         when "1111001100110" => index <= 8;
         when "1111001100111" => index <= 7;
         when "1111001101000" => index <= 9;
         when "1111001101001" => index <= 8;
         when "1111001101010" => index <= 8;
         when "1111001101011" => index <= 7;
         when "1111001101100" => index <= 8;
         when "1111001101101" => index <= 7;
         when "1111001101110" => index <= 8;
         when "1111001101111" => index <= 7;
         when "1111001110000" => index <= 9;
         when "1111001110001" => index <= 8;
         when "1111001110010" => index <= 8;
         when "1111001110011" => index <= 7;
         when "1111001110100" => index <= 8;
         when "1111001110101" => index <= 8;
         when "1111001110110" => index <= 8;
         when "1111001110111" => index <= 7;
         when "1111001111000" => index <= 8;
         when "1111001111001" => index <= 8;
         when "1111001111010" => index <= 8;
         when "1111001111011" => index <= 7;
         when "1111001111100" => index <= 8;
         when "1111001111101" => index <= 7;
         when "1111001111110" => index <= 7;
         when "1111001111111" => index <= 7;
         when "1111010000000" => index <= 11;
         when "1111010000001" => index <= 9;
         when "1111010000010" => index <= 9;
         when "1111010000011" => index <= 8;
         when "1111010000100" => index <= 10;
         when "1111010000101" => index <= 8;
         when "1111010000110" => index <= 8;
         when "1111010000111" => index <= 8;
         when "1111010001000" => index <= 10;
         when "1111010001001" => index <= 8;
         when "1111010001010" => index <= 9;
         when "1111010001011" => index <= 8;
         when "1111010001100" => index <= 9;
         when "1111010001101" => index <= 8;
         when "1111010001110" => index <= 8;
         when "1111010001111" => index <= 7;
         when "1111010010000" => index <= 10;
         when "1111010010001" => index <= 9;
         when "1111010010010" => index <= 9;
         when "1111010010011" => index <= 8;
         when "1111010010100" => index <= 9;
         when "1111010010101" => index <= 8;
         when "1111010010110" => index <= 8;
         when "1111010010111" => index <= 7;
         when "1111010011000" => index <= 9;
         when "1111010011001" => index <= 8;
         when "1111010011010" => index <= 8;
         when "1111010011011" => index <= 7;
         when "1111010011100" => index <= 8;
         when "1111010011101" => index <= 7;
         when "1111010011110" => index <= 8;
         when "1111010011111" => index <= 7;
         when "1111010100000" => index <= 10;
         when "1111010100001" => index <= 9;
         when "1111010100010" => index <= 9;
         when "1111010100011" => index <= 8;
         when "1111010100100" => index <= 9;
         when "1111010100101" => index <= 8;
         when "1111010100110" => index <= 8;
         when "1111010100111" => index <= 7;
         when "1111010101000" => index <= 9;
         when "1111010101001" => index <= 8;
         when "1111010101010" => index <= 8;
         when "1111010101011" => index <= 7;
         when "1111010101100" => index <= 8;
         when "1111010101101" => index <= 8;
         when "1111010101110" => index <= 8;
         when "1111010101111" => index <= 7;
         when "1111010110000" => index <= 9;
         when "1111010110001" => index <= 8;
         when "1111010110010" => index <= 8;
         when "1111010110011" => index <= 8;
         when "1111010110100" => index <= 8;
         when "1111010110101" => index <= 8;
         when "1111010110110" => index <= 8;
         when "1111010110111" => index <= 7;
         when "1111010111000" => index <= 9;
         when "1111010111001" => index <= 8;
         when "1111010111010" => index <= 8;
         when "1111010111011" => index <= 7;
         when "1111010111100" => index <= 8;
         when "1111010111101" => index <= 7;
         when "1111010111110" => index <= 7;
         when "1111010111111" => index <= 7;
         when "1111011000000" => index <= 10;
         when "1111011000001" => index <= 9;
         when "1111011000010" => index <= 9;
         when "1111011000011" => index <= 8;
         when "1111011000100" => index <= 9;
         when "1111011000101" => index <= 8;
         when "1111011000110" => index <= 8;
         when "1111011000111" => index <= 7;
         when "1111011001000" => index <= 9;
         when "1111011001001" => index <= 8;
         when "1111011001010" => index <= 8;
         when "1111011001011" => index <= 8;
         when "1111011001100" => index <= 8;
         when "1111011001101" => index <= 8;
         when "1111011001110" => index <= 8;
         when "1111011001111" => index <= 7;
         when "1111011010000" => index <= 9;
         when "1111011010001" => index <= 8;
         when "1111011010010" => index <= 8;
         when "1111011010011" => index <= 8;
         when "1111011010100" => index <= 9;
         when "1111011010101" => index <= 8;
         when "1111011010110" => index <= 8;
         when "1111011010111" => index <= 7;
         when "1111011011000" => index <= 9;
         when "1111011011001" => index <= 8;
         when "1111011011010" => index <= 8;
         when "1111011011011" => index <= 7;
         when "1111011011100" => index <= 8;
         when "1111011011101" => index <= 7;
         when "1111011011110" => index <= 8;
         when "1111011011111" => index <= 7;
         when "1111011100000" => index <= 10;
         when "1111011100001" => index <= 8;
         when "1111011100010" => index <= 9;
         when "1111011100011" => index <= 8;
         when "1111011100100" => index <= 9;
         when "1111011100101" => index <= 8;
         when "1111011100110" => index <= 8;
         when "1111011100111" => index <= 7;
         when "1111011101000" => index <= 9;
         when "1111011101001" => index <= 8;
         when "1111011101010" => index <= 8;
         when "1111011101011" => index <= 7;
         when "1111011101100" => index <= 8;
         when "1111011101101" => index <= 8;
         when "1111011101110" => index <= 8;
         when "1111011101111" => index <= 7;
         when "1111011110000" => index <= 9;
         when "1111011110001" => index <= 8;
         when "1111011110010" => index <= 8;
         when "1111011110011" => index <= 8;
         when "1111011110100" => index <= 8;
         when "1111011110101" => index <= 8;
         when "1111011110110" => index <= 8;
         when "1111011110111" => index <= 7;
         when "1111011111000" => index <= 8;
         when "1111011111001" => index <= 8;
         when "1111011111010" => index <= 8;
         when "1111011111011" => index <= 7;
         when "1111011111100" => index <= 8;
         when "1111011111101" => index <= 7;
         when "1111011111110" => index <= 7;
         when "1111011111111" => index <= 7;
         when "1111100000000" => index <= 11;
         when "1111100000001" => index <= 9;
         when "1111100000010" => index <= 10;
         when "1111100000011" => index <= 8;
         when "1111100000100" => index <= 10;
         when "1111100000101" => index <= 8;
         when "1111100000110" => index <= 9;
         when "1111100000111" => index <= 8;
         when "1111100001000" => index <= 10;
         when "1111100001001" => index <= 9;
         when "1111100001010" => index <= 9;
         when "1111100001011" => index <= 8;
         when "1111100001100" => index <= 9;
         when "1111100001101" => index <= 8;
         when "1111100001110" => index <= 8;
         when "1111100001111" => index <= 7;
         when "1111100010000" => index <= 10;
         when "1111100010001" => index <= 9;
         when "1111100010010" => index <= 9;
         when "1111100010011" => index <= 8;
         when "1111100010100" => index <= 9;
         when "1111100010101" => index <= 8;
         when "1111100010110" => index <= 8;
         when "1111100010111" => index <= 7;
         when "1111100011000" => index <= 9;
         when "1111100011001" => index <= 8;
         when "1111100011010" => index <= 8;
         when "1111100011011" => index <= 7;
         when "1111100011100" => index <= 8;
         when "1111100011101" => index <= 8;
         when "1111100011110" => index <= 8;
         when "1111100011111" => index <= 7;
         when "1111100100000" => index <= 10;
         when "1111100100001" => index <= 9;
         when "1111100100010" => index <= 9;
         when "1111100100011" => index <= 8;
         when "1111100100100" => index <= 9;
         when "1111100100101" => index <= 8;
         when "1111100100110" => index <= 8;
         when "1111100100111" => index <= 7;
         when "1111100101000" => index <= 9;
         when "1111100101001" => index <= 8;
         when "1111100101010" => index <= 8;
         when "1111100101011" => index <= 8;
         when "1111100101100" => index <= 8;
         when "1111100101101" => index <= 8;
         when "1111100101110" => index <= 8;
         when "1111100101111" => index <= 7;
         when "1111100110000" => index <= 9;
         when "1111100110001" => index <= 8;
         when "1111100110010" => index <= 8;
         when "1111100110011" => index <= 8;
         when "1111100110100" => index <= 9;
         when "1111100110101" => index <= 8;
         when "1111100110110" => index <= 8;
         when "1111100110111" => index <= 7;
         when "1111100111000" => index <= 9;
         when "1111100111001" => index <= 8;
         when "1111100111010" => index <= 8;
         when "1111100111011" => index <= 7;
         when "1111100111100" => index <= 8;
         when "1111100111101" => index <= 7;
         when "1111100111110" => index <= 8;
         when "1111100111111" => index <= 7;
         when "1111101000000" => index <= 10;
         when "1111101000001" => index <= 9;
         when "1111101000010" => index <= 9;
         when "1111101000011" => index <= 8;
         when "1111101000100" => index <= 9;
         when "1111101000101" => index <= 8;
         when "1111101000110" => index <= 8;
         when "1111101000111" => index <= 8;
         when "1111101001000" => index <= 9;
         when "1111101001001" => index <= 8;
         when "1111101001010" => index <= 8;
         when "1111101001011" => index <= 8;
         when "1111101001100" => index <= 9;
         when "1111101001101" => index <= 8;
         when "1111101001110" => index <= 8;
         when "1111101001111" => index <= 7;
         when "1111101010000" => index <= 10;
         when "1111101010001" => index <= 8;
         when "1111101010010" => index <= 9;
         when "1111101010011" => index <= 8;
         when "1111101010100" => index <= 9;
         when "1111101010101" => index <= 8;
         when "1111101010110" => index <= 8;
         when "1111101010111" => index <= 7;
         when "1111101011000" => index <= 9;
         when "1111101011001" => index <= 8;
         when "1111101011010" => index <= 8;
         when "1111101011011" => index <= 7;
         when "1111101011100" => index <= 8;
         when "1111101011101" => index <= 8;
         when "1111101011110" => index <= 8;
         when "1111101011111" => index <= 7;
         when "1111101100000" => index <= 10;
         when "1111101100001" => index <= 9;
         when "1111101100010" => index <= 9;
         when "1111101100011" => index <= 8;
         when "1111101100100" => index <= 9;
         when "1111101100101" => index <= 8;
         when "1111101100110" => index <= 8;
         when "1111101100111" => index <= 7;
         when "1111101101000" => index <= 9;
         when "1111101101001" => index <= 8;
         when "1111101101010" => index <= 8;
         when "1111101101011" => index <= 8;
         when "1111101101100" => index <= 8;
         when "1111101101101" => index <= 8;
         when "1111101101110" => index <= 8;
         when "1111101101111" => index <= 7;
         when "1111101110000" => index <= 9;
         when "1111101110001" => index <= 8;
         when "1111101110010" => index <= 8;
         when "1111101110011" => index <= 8;
         when "1111101110100" => index <= 8;
         when "1111101110101" => index <= 8;
         when "1111101110110" => index <= 8;
         when "1111101110111" => index <= 7;
         when "1111101111000" => index <= 9;
         when "1111101111001" => index <= 8;
         when "1111101111010" => index <= 8;
         when "1111101111011" => index <= 7;
         when "1111101111100" => index <= 8;
         when "1111101111101" => index <= 7;
         when "1111101111110" => index <= 7;
         when "1111101111111" => index <= 7;
         when "1111110000000" => index <= 10;
         when "1111110000001" => index <= 9;
         when "1111110000010" => index <= 9;
         when "1111110000011" => index <= 8;
         when "1111110000100" => index <= 9;
         when "1111110000101" => index <= 8;
         when "1111110000110" => index <= 8;
         when "1111110000111" => index <= 8;
         when "1111110001000" => index <= 10;
         when "1111110001001" => index <= 8;
         when "1111110001010" => index <= 9;
         when "1111110001011" => index <= 8;
         when "1111110001100" => index <= 9;
         when "1111110001101" => index <= 8;
         when "1111110001110" => index <= 8;
         when "1111110001111" => index <= 7;
         when "1111110010000" => index <= 10;
         when "1111110010001" => index <= 9;
         when "1111110010010" => index <= 9;
         when "1111110010011" => index <= 8;
         when "1111110010100" => index <= 9;
         when "1111110010101" => index <= 8;
         when "1111110010110" => index <= 8;
         when "1111110010111" => index <= 7;
         when "1111110011000" => index <= 9;
         when "1111110011001" => index <= 8;
         when "1111110011010" => index <= 8;
         when "1111110011011" => index <= 8;
         when "1111110011100" => index <= 8;
         when "1111110011101" => index <= 8;
         when "1111110011110" => index <= 8;
         when "1111110011111" => index <= 7;
         when "1111110100000" => index <= 10;
         when "1111110100001" => index <= 9;
         when "1111110100010" => index <= 9;
         when "1111110100011" => index <= 8;
         when "1111110100100" => index <= 9;
         when "1111110100101" => index <= 8;
         when "1111110100110" => index <= 8;
         when "1111110100111" => index <= 8;
         when "1111110101000" => index <= 9;
         when "1111110101001" => index <= 8;
         when "1111110101010" => index <= 8;
         when "1111110101011" => index <= 8;
         when "1111110101100" => index <= 8;
         when "1111110101101" => index <= 8;
         when "1111110101110" => index <= 8;
         when "1111110101111" => index <= 7;
         when "1111110110000" => index <= 9;
         when "1111110110001" => index <= 8;
         when "1111110110010" => index <= 8;
         when "1111110110011" => index <= 8;
         when "1111110110100" => index <= 9;
         when "1111110110101" => index <= 8;
         when "1111110110110" => index <= 8;
         when "1111110110111" => index <= 7;
         when "1111110111000" => index <= 9;
         when "1111110111001" => index <= 8;
         when "1111110111010" => index <= 8;
         when "1111110111011" => index <= 7;
         when "1111110111100" => index <= 8;
         when "1111110111101" => index <= 7;
         when "1111110111110" => index <= 8;
         when "1111110111111" => index <= 7;
         when "1111111000000" => index <= 10;
         when "1111111000001" => index <= 9;
         when "1111111000010" => index <= 9;
         when "1111111000011" => index <= 8;
         when "1111111000100" => index <= 9;
         when "1111111000101" => index <= 8;
         when "1111111000110" => index <= 8;
         when "1111111000111" => index <= 8;
         when "1111111001000" => index <= 9;
         when "1111111001001" => index <= 8;
         when "1111111001010" => index <= 8;
         when "1111111001011" => index <= 8;
         when "1111111001100" => index <= 9;
         when "1111111001101" => index <= 8;
         when "1111111001110" => index <= 8;
         when "1111111001111" => index <= 7;
         when "1111111010000" => index <= 9;
         when "1111111010001" => index <= 8;
         when "1111111010010" => index <= 9;
         when "1111111010011" => index <= 8;
         when "1111111010100" => index <= 9;
         when "1111111010101" => index <= 8;
         when "1111111010110" => index <= 8;
         when "1111111010111" => index <= 7;
         when "1111111011000" => index <= 9;
         when "1111111011001" => index <= 8;
         when "1111111011010" => index <= 8;
         when "1111111011011" => index <= 7;
         when "1111111011100" => index <= 8;
         when "1111111011101" => index <= 8;
         when "1111111011110" => index <= 8;
         when "1111111011111" => index <= 7;
         when "1111111100000" => index <= 10;
         when "1111111100001" => index <= 9;
         when "1111111100010" => index <= 9;
         when "1111111100011" => index <= 8;
         when "1111111100100" => index <= 9;
         when "1111111100101" => index <= 8;
         when "1111111100110" => index <= 8;
         when "1111111100111" => index <= 7;
         when "1111111101000" => index <= 9;
         when "1111111101001" => index <= 8;
         when "1111111101010" => index <= 8;
         when "1111111101011" => index <= 8;
         when "1111111101100" => index <= 8;
         when "1111111101101" => index <= 8;
         when "1111111101110" => index <= 8;
         when "1111111101111" => index <= 7;
         when "1111111110000" => index <= 9;
         when "1111111110001" => index <= 8;
         when "1111111110010" => index <= 8;
         when "1111111110011" => index <= 8;
         when "1111111110100" => index <= 8;
         when "1111111110101" => index <= 8;
         when "1111111110110" => index <= 8;
         when "1111111110111" => index <= 7;
         when "1111111111000" => index <= 8;
         when "1111111111001" => index <= 8;
         when "1111111111010" => index <= 8;
         when "1111111111011" => index <= 7;
         when "1111111111100" => index <= 8;
         when "1111111111101" => index <= 7;
         when "1111111111110" => index <= 8;
         when "1111111111111" => index <= 7;
         when others => index <= 0;
        end case;
      end if;
    end process;
  dout <= to_unsigned(index, NBITS);
  end generate;




end behavioral;
