library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

package bitonic_sort_pkg is
  type t_slm is array(natural range <>, natural range <>) of std_logic;
end package bitonic_sort_pkg;
